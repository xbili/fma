module fma_8x8(out_0, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15);
input [7:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15;
output [21:0] out_0;
wire [1897:0] wires;
assign wires[0] = in_0[0];
assign wires[1] = in_0[1];
assign wires[2] = in_0[2];
assign wires[3] = in_0[3];
assign wires[4] = in_0[4];
assign wires[5] = in_0[5];
assign wires[6] = in_0[6];
assign wires[7] = in_0[7];
assign wires[8] = in_1[0];
assign wires[9] = in_1[1];
assign wires[10] = in_1[2];
assign wires[11] = in_1[3];
assign wires[12] = in_1[4];
assign wires[13] = in_1[5];
assign wires[14] = in_1[6];
assign wires[15] = in_1[7];
assign wires[96] = in_2[0];
assign wires[97] = in_2[1];
assign wires[98] = in_2[2];
assign wires[99] = in_2[3];
assign wires[100] = in_2[4];
assign wires[101] = in_2[5];
assign wires[102] = in_2[6];
assign wires[103] = in_2[7];
assign wires[104] = in_3[0];
assign wires[105] = in_3[1];
assign wires[106] = in_3[2];
assign wires[107] = in_3[3];
assign wires[108] = in_3[4];
assign wires[109] = in_3[5];
assign wires[110] = in_3[6];
assign wires[111] = in_3[7];
assign wires[192] = in_4[0];
assign wires[193] = in_4[1];
assign wires[194] = in_4[2];
assign wires[195] = in_4[3];
assign wires[196] = in_4[4];
assign wires[197] = in_4[5];
assign wires[198] = in_4[6];
assign wires[199] = in_4[7];
assign wires[200] = in_5[0];
assign wires[201] = in_5[1];
assign wires[202] = in_5[2];
assign wires[203] = in_5[3];
assign wires[204] = in_5[4];
assign wires[205] = in_5[5];
assign wires[206] = in_5[6];
assign wires[207] = in_5[7];
assign wires[288] = in_6[0];
assign wires[289] = in_6[1];
assign wires[290] = in_6[2];
assign wires[291] = in_6[3];
assign wires[292] = in_6[4];
assign wires[293] = in_6[5];
assign wires[294] = in_6[6];
assign wires[295] = in_6[7];
assign wires[296] = in_7[0];
assign wires[297] = in_7[1];
assign wires[298] = in_7[2];
assign wires[299] = in_7[3];
assign wires[300] = in_7[4];
assign wires[301] = in_7[5];
assign wires[302] = in_7[6];
assign wires[303] = in_7[7];
assign wires[384] = in_8[0];
assign wires[385] = in_8[1];
assign wires[386] = in_8[2];
assign wires[387] = in_8[3];
assign wires[388] = in_8[4];
assign wires[389] = in_8[5];
assign wires[390] = in_8[6];
assign wires[391] = in_8[7];
assign wires[392] = in_9[0];
assign wires[393] = in_9[1];
assign wires[394] = in_9[2];
assign wires[395] = in_9[3];
assign wires[396] = in_9[4];
assign wires[397] = in_9[5];
assign wires[398] = in_9[6];
assign wires[399] = in_9[7];
assign wires[480] = in_10[0];
assign wires[481] = in_10[1];
assign wires[482] = in_10[2];
assign wires[483] = in_10[3];
assign wires[484] = in_10[4];
assign wires[485] = in_10[5];
assign wires[486] = in_10[6];
assign wires[487] = in_10[7];
assign wires[488] = in_11[0];
assign wires[489] = in_11[1];
assign wires[490] = in_11[2];
assign wires[491] = in_11[3];
assign wires[492] = in_11[4];
assign wires[493] = in_11[5];
assign wires[494] = in_11[6];
assign wires[495] = in_11[7];
assign wires[576] = in_12[0];
assign wires[577] = in_12[1];
assign wires[578] = in_12[2];
assign wires[579] = in_12[3];
assign wires[580] = in_12[4];
assign wires[581] = in_12[5];
assign wires[582] = in_12[6];
assign wires[583] = in_12[7];
assign wires[584] = in_13[0];
assign wires[585] = in_13[1];
assign wires[586] = in_13[2];
assign wires[587] = in_13[3];
assign wires[588] = in_13[4];
assign wires[589] = in_13[5];
assign wires[590] = in_13[6];
assign wires[591] = in_13[7];
assign wires[672] = in_14[0];
assign wires[673] = in_14[1];
assign wires[674] = in_14[2];
assign wires[675] = in_14[3];
assign wires[676] = in_14[4];
assign wires[677] = in_14[5];
assign wires[678] = in_14[6];
assign wires[679] = in_14[7];
assign wires[680] = in_15[0];
assign wires[681] = in_15[1];
assign wires[682] = in_15[2];
assign wires[683] = in_15[3];
assign wires[684] = in_15[4];
assign wires[685] = in_15[5];
assign wires[686] = in_15[6];
assign wires[687] = in_15[7];
assign out_0[0] = wires[1120];
assign out_0[1] = wires[1522];
assign out_0[2] = wires[1634];
assign out_0[3] = wires[1712];
assign out_0[4] = wires[1770];
assign out_0[5] = wires[1812];
assign out_0[6] = wires[1842];
assign out_0[7] = wires[1870];
assign out_0[8] = wires[1872];
assign out_0[9] = wires[1874];
assign out_0[10] = wires[1876];
assign out_0[11] = wires[1878];
assign out_0[12] = wires[1880];
assign out_0[13] = wires[1882];
assign out_0[14] = wires[1884];
assign out_0[15] = wires[1886];
assign out_0[16] = wires[1888];
assign out_0[17] = wires[1890];
assign out_0[18] = wires[1892];
assign out_0[19] = wires[1894];
assign out_0[20] = wires[1896];
assign out_0[21] = wires[1897];
and(wires[16], wires[8], wires[0]);
and(wires[17], wires[9], wires[0]);
and(wires[18], wires[10], wires[0]);
and(wires[19], wires[11], wires[0]);
and(wires[20], wires[12], wires[0]);
and(wires[21], wires[13], wires[0]);
and(wires[22], wires[14], wires[0]);
and(wires[23], wires[15], wires[0]);
not(wires[24], wires[23]);
and(wires[25], wires[8], wires[1]);
and(wires[26], wires[9], wires[1]);
and(wires[27], wires[10], wires[1]);
and(wires[28], wires[11], wires[1]);
and(wires[29], wires[12], wires[1]);
and(wires[30], wires[13], wires[1]);
and(wires[31], wires[14], wires[1]);
and(wires[32], wires[15], wires[1]);
not(wires[33], wires[32]);
and(wires[34], wires[8], wires[2]);
and(wires[35], wires[9], wires[2]);
and(wires[36], wires[10], wires[2]);
and(wires[37], wires[11], wires[2]);
and(wires[38], wires[12], wires[2]);
and(wires[39], wires[13], wires[2]);
and(wires[40], wires[14], wires[2]);
and(wires[41], wires[15], wires[2]);
not(wires[42], wires[41]);
and(wires[43], wires[8], wires[3]);
and(wires[44], wires[9], wires[3]);
and(wires[45], wires[10], wires[3]);
and(wires[46], wires[11], wires[3]);
and(wires[47], wires[12], wires[3]);
and(wires[48], wires[13], wires[3]);
and(wires[49], wires[14], wires[3]);
and(wires[50], wires[15], wires[3]);
not(wires[51], wires[50]);
and(wires[52], wires[8], wires[4]);
and(wires[53], wires[9], wires[4]);
and(wires[54], wires[10], wires[4]);
and(wires[55], wires[11], wires[4]);
and(wires[56], wires[12], wires[4]);
and(wires[57], wires[13], wires[4]);
and(wires[58], wires[14], wires[4]);
and(wires[59], wires[15], wires[4]);
not(wires[60], wires[59]);
and(wires[61], wires[8], wires[5]);
and(wires[62], wires[9], wires[5]);
and(wires[63], wires[10], wires[5]);
and(wires[64], wires[11], wires[5]);
and(wires[65], wires[12], wires[5]);
and(wires[66], wires[13], wires[5]);
and(wires[67], wires[14], wires[5]);
and(wires[68], wires[15], wires[5]);
not(wires[69], wires[68]);
and(wires[70], wires[8], wires[6]);
and(wires[71], wires[9], wires[6]);
and(wires[72], wires[10], wires[6]);
and(wires[73], wires[11], wires[6]);
and(wires[74], wires[12], wires[6]);
and(wires[75], wires[13], wires[6]);
and(wires[76], wires[14], wires[6]);
and(wires[77], wires[15], wires[6]);
not(wires[78], wires[77]);
and(wires[80], wires[8], wires[7]);
not(wires[81], wires[80]);
and(wires[82], wires[9], wires[7]);
not(wires[83], wires[82]);
and(wires[84], wires[10], wires[7]);
not(wires[85], wires[84]);
and(wires[86], wires[11], wires[7]);
not(wires[87], wires[86]);
and(wires[88], wires[12], wires[7]);
not(wires[89], wires[88]);
and(wires[90], wires[13], wires[7]);
not(wires[91], wires[90]);
and(wires[92], wires[14], wires[7]);
not(wires[93], wires[92]);
and(wires[94], wires[15], wires[7]);
and(wires[112], wires[104], wires[96]);
and(wires[113], wires[105], wires[96]);
and(wires[114], wires[106], wires[96]);
and(wires[115], wires[107], wires[96]);
and(wires[116], wires[108], wires[96]);
and(wires[117], wires[109], wires[96]);
and(wires[118], wires[110], wires[96]);
and(wires[119], wires[111], wires[96]);
not(wires[120], wires[119]);
and(wires[121], wires[104], wires[97]);
and(wires[122], wires[105], wires[97]);
and(wires[123], wires[106], wires[97]);
and(wires[124], wires[107], wires[97]);
and(wires[125], wires[108], wires[97]);
and(wires[126], wires[109], wires[97]);
and(wires[127], wires[110], wires[97]);
and(wires[128], wires[111], wires[97]);
not(wires[129], wires[128]);
and(wires[130], wires[104], wires[98]);
and(wires[131], wires[105], wires[98]);
and(wires[132], wires[106], wires[98]);
and(wires[133], wires[107], wires[98]);
and(wires[134], wires[108], wires[98]);
and(wires[135], wires[109], wires[98]);
and(wires[136], wires[110], wires[98]);
and(wires[137], wires[111], wires[98]);
not(wires[138], wires[137]);
and(wires[139], wires[104], wires[99]);
and(wires[140], wires[105], wires[99]);
and(wires[141], wires[106], wires[99]);
and(wires[142], wires[107], wires[99]);
and(wires[143], wires[108], wires[99]);
and(wires[144], wires[109], wires[99]);
and(wires[145], wires[110], wires[99]);
and(wires[146], wires[111], wires[99]);
not(wires[147], wires[146]);
and(wires[148], wires[104], wires[100]);
and(wires[149], wires[105], wires[100]);
and(wires[150], wires[106], wires[100]);
and(wires[151], wires[107], wires[100]);
and(wires[152], wires[108], wires[100]);
and(wires[153], wires[109], wires[100]);
and(wires[154], wires[110], wires[100]);
and(wires[155], wires[111], wires[100]);
not(wires[156], wires[155]);
and(wires[157], wires[104], wires[101]);
and(wires[158], wires[105], wires[101]);
and(wires[159], wires[106], wires[101]);
and(wires[160], wires[107], wires[101]);
and(wires[161], wires[108], wires[101]);
and(wires[162], wires[109], wires[101]);
and(wires[163], wires[110], wires[101]);
and(wires[164], wires[111], wires[101]);
not(wires[165], wires[164]);
and(wires[166], wires[104], wires[102]);
and(wires[167], wires[105], wires[102]);
and(wires[168], wires[106], wires[102]);
and(wires[169], wires[107], wires[102]);
and(wires[170], wires[108], wires[102]);
and(wires[171], wires[109], wires[102]);
and(wires[172], wires[110], wires[102]);
and(wires[173], wires[111], wires[102]);
not(wires[174], wires[173]);
and(wires[176], wires[104], wires[103]);
not(wires[177], wires[176]);
and(wires[178], wires[105], wires[103]);
not(wires[179], wires[178]);
and(wires[180], wires[106], wires[103]);
not(wires[181], wires[180]);
and(wires[182], wires[107], wires[103]);
not(wires[183], wires[182]);
and(wires[184], wires[108], wires[103]);
not(wires[185], wires[184]);
and(wires[186], wires[109], wires[103]);
not(wires[187], wires[186]);
and(wires[188], wires[110], wires[103]);
not(wires[189], wires[188]);
and(wires[190], wires[111], wires[103]);
and(wires[208], wires[200], wires[192]);
and(wires[209], wires[201], wires[192]);
and(wires[210], wires[202], wires[192]);
and(wires[211], wires[203], wires[192]);
and(wires[212], wires[204], wires[192]);
and(wires[213], wires[205], wires[192]);
and(wires[214], wires[206], wires[192]);
and(wires[215], wires[207], wires[192]);
not(wires[216], wires[215]);
and(wires[217], wires[200], wires[193]);
and(wires[218], wires[201], wires[193]);
and(wires[219], wires[202], wires[193]);
and(wires[220], wires[203], wires[193]);
and(wires[221], wires[204], wires[193]);
and(wires[222], wires[205], wires[193]);
and(wires[223], wires[206], wires[193]);
and(wires[224], wires[207], wires[193]);
not(wires[225], wires[224]);
and(wires[226], wires[200], wires[194]);
and(wires[227], wires[201], wires[194]);
and(wires[228], wires[202], wires[194]);
and(wires[229], wires[203], wires[194]);
and(wires[230], wires[204], wires[194]);
and(wires[231], wires[205], wires[194]);
and(wires[232], wires[206], wires[194]);
and(wires[233], wires[207], wires[194]);
not(wires[234], wires[233]);
and(wires[235], wires[200], wires[195]);
and(wires[236], wires[201], wires[195]);
and(wires[237], wires[202], wires[195]);
and(wires[238], wires[203], wires[195]);
and(wires[239], wires[204], wires[195]);
and(wires[240], wires[205], wires[195]);
and(wires[241], wires[206], wires[195]);
and(wires[242], wires[207], wires[195]);
not(wires[243], wires[242]);
and(wires[244], wires[200], wires[196]);
and(wires[245], wires[201], wires[196]);
and(wires[246], wires[202], wires[196]);
and(wires[247], wires[203], wires[196]);
and(wires[248], wires[204], wires[196]);
and(wires[249], wires[205], wires[196]);
and(wires[250], wires[206], wires[196]);
and(wires[251], wires[207], wires[196]);
not(wires[252], wires[251]);
and(wires[253], wires[200], wires[197]);
and(wires[254], wires[201], wires[197]);
and(wires[255], wires[202], wires[197]);
and(wires[256], wires[203], wires[197]);
and(wires[257], wires[204], wires[197]);
and(wires[258], wires[205], wires[197]);
and(wires[259], wires[206], wires[197]);
and(wires[260], wires[207], wires[197]);
not(wires[261], wires[260]);
and(wires[262], wires[200], wires[198]);
and(wires[263], wires[201], wires[198]);
and(wires[264], wires[202], wires[198]);
and(wires[265], wires[203], wires[198]);
and(wires[266], wires[204], wires[198]);
and(wires[267], wires[205], wires[198]);
and(wires[268], wires[206], wires[198]);
and(wires[269], wires[207], wires[198]);
not(wires[270], wires[269]);
and(wires[272], wires[200], wires[199]);
not(wires[273], wires[272]);
and(wires[274], wires[201], wires[199]);
not(wires[275], wires[274]);
and(wires[276], wires[202], wires[199]);
not(wires[277], wires[276]);
and(wires[278], wires[203], wires[199]);
not(wires[279], wires[278]);
and(wires[280], wires[204], wires[199]);
not(wires[281], wires[280]);
and(wires[282], wires[205], wires[199]);
not(wires[283], wires[282]);
and(wires[284], wires[206], wires[199]);
not(wires[285], wires[284]);
and(wires[286], wires[207], wires[199]);
and(wires[304], wires[296], wires[288]);
and(wires[305], wires[297], wires[288]);
and(wires[306], wires[298], wires[288]);
and(wires[307], wires[299], wires[288]);
and(wires[308], wires[300], wires[288]);
and(wires[309], wires[301], wires[288]);
and(wires[310], wires[302], wires[288]);
and(wires[311], wires[303], wires[288]);
not(wires[312], wires[311]);
and(wires[313], wires[296], wires[289]);
and(wires[314], wires[297], wires[289]);
and(wires[315], wires[298], wires[289]);
and(wires[316], wires[299], wires[289]);
and(wires[317], wires[300], wires[289]);
and(wires[318], wires[301], wires[289]);
and(wires[319], wires[302], wires[289]);
and(wires[320], wires[303], wires[289]);
not(wires[321], wires[320]);
and(wires[322], wires[296], wires[290]);
and(wires[323], wires[297], wires[290]);
and(wires[324], wires[298], wires[290]);
and(wires[325], wires[299], wires[290]);
and(wires[326], wires[300], wires[290]);
and(wires[327], wires[301], wires[290]);
and(wires[328], wires[302], wires[290]);
and(wires[329], wires[303], wires[290]);
not(wires[330], wires[329]);
and(wires[331], wires[296], wires[291]);
and(wires[332], wires[297], wires[291]);
and(wires[333], wires[298], wires[291]);
and(wires[334], wires[299], wires[291]);
and(wires[335], wires[300], wires[291]);
and(wires[336], wires[301], wires[291]);
and(wires[337], wires[302], wires[291]);
and(wires[338], wires[303], wires[291]);
not(wires[339], wires[338]);
and(wires[340], wires[296], wires[292]);
and(wires[341], wires[297], wires[292]);
and(wires[342], wires[298], wires[292]);
and(wires[343], wires[299], wires[292]);
and(wires[344], wires[300], wires[292]);
and(wires[345], wires[301], wires[292]);
and(wires[346], wires[302], wires[292]);
and(wires[347], wires[303], wires[292]);
not(wires[348], wires[347]);
and(wires[349], wires[296], wires[293]);
and(wires[350], wires[297], wires[293]);
and(wires[351], wires[298], wires[293]);
and(wires[352], wires[299], wires[293]);
and(wires[353], wires[300], wires[293]);
and(wires[354], wires[301], wires[293]);
and(wires[355], wires[302], wires[293]);
and(wires[356], wires[303], wires[293]);
not(wires[357], wires[356]);
and(wires[358], wires[296], wires[294]);
and(wires[359], wires[297], wires[294]);
and(wires[360], wires[298], wires[294]);
and(wires[361], wires[299], wires[294]);
and(wires[362], wires[300], wires[294]);
and(wires[363], wires[301], wires[294]);
and(wires[364], wires[302], wires[294]);
and(wires[365], wires[303], wires[294]);
not(wires[366], wires[365]);
and(wires[368], wires[296], wires[295]);
not(wires[369], wires[368]);
and(wires[370], wires[297], wires[295]);
not(wires[371], wires[370]);
and(wires[372], wires[298], wires[295]);
not(wires[373], wires[372]);
and(wires[374], wires[299], wires[295]);
not(wires[375], wires[374]);
and(wires[376], wires[300], wires[295]);
not(wires[377], wires[376]);
and(wires[378], wires[301], wires[295]);
not(wires[379], wires[378]);
and(wires[380], wires[302], wires[295]);
not(wires[381], wires[380]);
and(wires[382], wires[303], wires[295]);
and(wires[400], wires[392], wires[384]);
and(wires[401], wires[393], wires[384]);
and(wires[402], wires[394], wires[384]);
and(wires[403], wires[395], wires[384]);
and(wires[404], wires[396], wires[384]);
and(wires[405], wires[397], wires[384]);
and(wires[406], wires[398], wires[384]);
and(wires[407], wires[399], wires[384]);
not(wires[408], wires[407]);
and(wires[409], wires[392], wires[385]);
and(wires[410], wires[393], wires[385]);
and(wires[411], wires[394], wires[385]);
and(wires[412], wires[395], wires[385]);
and(wires[413], wires[396], wires[385]);
and(wires[414], wires[397], wires[385]);
and(wires[415], wires[398], wires[385]);
and(wires[416], wires[399], wires[385]);
not(wires[417], wires[416]);
and(wires[418], wires[392], wires[386]);
and(wires[419], wires[393], wires[386]);
and(wires[420], wires[394], wires[386]);
and(wires[421], wires[395], wires[386]);
and(wires[422], wires[396], wires[386]);
and(wires[423], wires[397], wires[386]);
and(wires[424], wires[398], wires[386]);
and(wires[425], wires[399], wires[386]);
not(wires[426], wires[425]);
and(wires[427], wires[392], wires[387]);
and(wires[428], wires[393], wires[387]);
and(wires[429], wires[394], wires[387]);
and(wires[430], wires[395], wires[387]);
and(wires[431], wires[396], wires[387]);
and(wires[432], wires[397], wires[387]);
and(wires[433], wires[398], wires[387]);
and(wires[434], wires[399], wires[387]);
not(wires[435], wires[434]);
and(wires[436], wires[392], wires[388]);
and(wires[437], wires[393], wires[388]);
and(wires[438], wires[394], wires[388]);
and(wires[439], wires[395], wires[388]);
and(wires[440], wires[396], wires[388]);
and(wires[441], wires[397], wires[388]);
and(wires[442], wires[398], wires[388]);
and(wires[443], wires[399], wires[388]);
not(wires[444], wires[443]);
and(wires[445], wires[392], wires[389]);
and(wires[446], wires[393], wires[389]);
and(wires[447], wires[394], wires[389]);
and(wires[448], wires[395], wires[389]);
and(wires[449], wires[396], wires[389]);
and(wires[450], wires[397], wires[389]);
and(wires[451], wires[398], wires[389]);
and(wires[452], wires[399], wires[389]);
not(wires[453], wires[452]);
and(wires[454], wires[392], wires[390]);
and(wires[455], wires[393], wires[390]);
and(wires[456], wires[394], wires[390]);
and(wires[457], wires[395], wires[390]);
and(wires[458], wires[396], wires[390]);
and(wires[459], wires[397], wires[390]);
and(wires[460], wires[398], wires[390]);
and(wires[461], wires[399], wires[390]);
not(wires[462], wires[461]);
and(wires[464], wires[392], wires[391]);
not(wires[465], wires[464]);
and(wires[466], wires[393], wires[391]);
not(wires[467], wires[466]);
and(wires[468], wires[394], wires[391]);
not(wires[469], wires[468]);
and(wires[470], wires[395], wires[391]);
not(wires[471], wires[470]);
and(wires[472], wires[396], wires[391]);
not(wires[473], wires[472]);
and(wires[474], wires[397], wires[391]);
not(wires[475], wires[474]);
and(wires[476], wires[398], wires[391]);
not(wires[477], wires[476]);
and(wires[478], wires[399], wires[391]);
and(wires[496], wires[488], wires[480]);
and(wires[497], wires[489], wires[480]);
and(wires[498], wires[490], wires[480]);
and(wires[499], wires[491], wires[480]);
and(wires[500], wires[492], wires[480]);
and(wires[501], wires[493], wires[480]);
and(wires[502], wires[494], wires[480]);
and(wires[503], wires[495], wires[480]);
not(wires[504], wires[503]);
and(wires[505], wires[488], wires[481]);
and(wires[506], wires[489], wires[481]);
and(wires[507], wires[490], wires[481]);
and(wires[508], wires[491], wires[481]);
and(wires[509], wires[492], wires[481]);
and(wires[510], wires[493], wires[481]);
and(wires[511], wires[494], wires[481]);
and(wires[512], wires[495], wires[481]);
not(wires[513], wires[512]);
and(wires[514], wires[488], wires[482]);
and(wires[515], wires[489], wires[482]);
and(wires[516], wires[490], wires[482]);
and(wires[517], wires[491], wires[482]);
and(wires[518], wires[492], wires[482]);
and(wires[519], wires[493], wires[482]);
and(wires[520], wires[494], wires[482]);
and(wires[521], wires[495], wires[482]);
not(wires[522], wires[521]);
and(wires[523], wires[488], wires[483]);
and(wires[524], wires[489], wires[483]);
and(wires[525], wires[490], wires[483]);
and(wires[526], wires[491], wires[483]);
and(wires[527], wires[492], wires[483]);
and(wires[528], wires[493], wires[483]);
and(wires[529], wires[494], wires[483]);
and(wires[530], wires[495], wires[483]);
not(wires[531], wires[530]);
and(wires[532], wires[488], wires[484]);
and(wires[533], wires[489], wires[484]);
and(wires[534], wires[490], wires[484]);
and(wires[535], wires[491], wires[484]);
and(wires[536], wires[492], wires[484]);
and(wires[537], wires[493], wires[484]);
and(wires[538], wires[494], wires[484]);
and(wires[539], wires[495], wires[484]);
not(wires[540], wires[539]);
and(wires[541], wires[488], wires[485]);
and(wires[542], wires[489], wires[485]);
and(wires[543], wires[490], wires[485]);
and(wires[544], wires[491], wires[485]);
and(wires[545], wires[492], wires[485]);
and(wires[546], wires[493], wires[485]);
and(wires[547], wires[494], wires[485]);
and(wires[548], wires[495], wires[485]);
not(wires[549], wires[548]);
and(wires[550], wires[488], wires[486]);
and(wires[551], wires[489], wires[486]);
and(wires[552], wires[490], wires[486]);
and(wires[553], wires[491], wires[486]);
and(wires[554], wires[492], wires[486]);
and(wires[555], wires[493], wires[486]);
and(wires[556], wires[494], wires[486]);
and(wires[557], wires[495], wires[486]);
not(wires[558], wires[557]);
and(wires[560], wires[488], wires[487]);
not(wires[561], wires[560]);
and(wires[562], wires[489], wires[487]);
not(wires[563], wires[562]);
and(wires[564], wires[490], wires[487]);
not(wires[565], wires[564]);
and(wires[566], wires[491], wires[487]);
not(wires[567], wires[566]);
and(wires[568], wires[492], wires[487]);
not(wires[569], wires[568]);
and(wires[570], wires[493], wires[487]);
not(wires[571], wires[570]);
and(wires[572], wires[494], wires[487]);
not(wires[573], wires[572]);
and(wires[574], wires[495], wires[487]);
and(wires[592], wires[584], wires[576]);
and(wires[593], wires[585], wires[576]);
and(wires[594], wires[586], wires[576]);
and(wires[595], wires[587], wires[576]);
and(wires[596], wires[588], wires[576]);
and(wires[597], wires[589], wires[576]);
and(wires[598], wires[590], wires[576]);
and(wires[599], wires[591], wires[576]);
not(wires[600], wires[599]);
and(wires[601], wires[584], wires[577]);
and(wires[602], wires[585], wires[577]);
and(wires[603], wires[586], wires[577]);
and(wires[604], wires[587], wires[577]);
and(wires[605], wires[588], wires[577]);
and(wires[606], wires[589], wires[577]);
and(wires[607], wires[590], wires[577]);
and(wires[608], wires[591], wires[577]);
not(wires[609], wires[608]);
and(wires[610], wires[584], wires[578]);
and(wires[611], wires[585], wires[578]);
and(wires[612], wires[586], wires[578]);
and(wires[613], wires[587], wires[578]);
and(wires[614], wires[588], wires[578]);
and(wires[615], wires[589], wires[578]);
and(wires[616], wires[590], wires[578]);
and(wires[617], wires[591], wires[578]);
not(wires[618], wires[617]);
and(wires[619], wires[584], wires[579]);
and(wires[620], wires[585], wires[579]);
and(wires[621], wires[586], wires[579]);
and(wires[622], wires[587], wires[579]);
and(wires[623], wires[588], wires[579]);
and(wires[624], wires[589], wires[579]);
and(wires[625], wires[590], wires[579]);
and(wires[626], wires[591], wires[579]);
not(wires[627], wires[626]);
and(wires[628], wires[584], wires[580]);
and(wires[629], wires[585], wires[580]);
and(wires[630], wires[586], wires[580]);
and(wires[631], wires[587], wires[580]);
and(wires[632], wires[588], wires[580]);
and(wires[633], wires[589], wires[580]);
and(wires[634], wires[590], wires[580]);
and(wires[635], wires[591], wires[580]);
not(wires[636], wires[635]);
and(wires[637], wires[584], wires[581]);
and(wires[638], wires[585], wires[581]);
and(wires[639], wires[586], wires[581]);
and(wires[640], wires[587], wires[581]);
and(wires[641], wires[588], wires[581]);
and(wires[642], wires[589], wires[581]);
and(wires[643], wires[590], wires[581]);
and(wires[644], wires[591], wires[581]);
not(wires[645], wires[644]);
and(wires[646], wires[584], wires[582]);
and(wires[647], wires[585], wires[582]);
and(wires[648], wires[586], wires[582]);
and(wires[649], wires[587], wires[582]);
and(wires[650], wires[588], wires[582]);
and(wires[651], wires[589], wires[582]);
and(wires[652], wires[590], wires[582]);
and(wires[653], wires[591], wires[582]);
not(wires[654], wires[653]);
and(wires[656], wires[584], wires[583]);
not(wires[657], wires[656]);
and(wires[658], wires[585], wires[583]);
not(wires[659], wires[658]);
and(wires[660], wires[586], wires[583]);
not(wires[661], wires[660]);
and(wires[662], wires[587], wires[583]);
not(wires[663], wires[662]);
and(wires[664], wires[588], wires[583]);
not(wires[665], wires[664]);
and(wires[666], wires[589], wires[583]);
not(wires[667], wires[666]);
and(wires[668], wires[590], wires[583]);
not(wires[669], wires[668]);
and(wires[670], wires[591], wires[583]);
and(wires[688], wires[680], wires[672]);
and(wires[689], wires[681], wires[672]);
and(wires[690], wires[682], wires[672]);
and(wires[691], wires[683], wires[672]);
and(wires[692], wires[684], wires[672]);
and(wires[693], wires[685], wires[672]);
and(wires[694], wires[686], wires[672]);
and(wires[695], wires[687], wires[672]);
not(wires[696], wires[695]);
and(wires[697], wires[680], wires[673]);
and(wires[698], wires[681], wires[673]);
and(wires[699], wires[682], wires[673]);
and(wires[700], wires[683], wires[673]);
and(wires[701], wires[684], wires[673]);
and(wires[702], wires[685], wires[673]);
and(wires[703], wires[686], wires[673]);
and(wires[704], wires[687], wires[673]);
not(wires[705], wires[704]);
and(wires[706], wires[680], wires[674]);
and(wires[707], wires[681], wires[674]);
and(wires[708], wires[682], wires[674]);
and(wires[709], wires[683], wires[674]);
and(wires[710], wires[684], wires[674]);
and(wires[711], wires[685], wires[674]);
and(wires[712], wires[686], wires[674]);
and(wires[713], wires[687], wires[674]);
not(wires[714], wires[713]);
and(wires[715], wires[680], wires[675]);
and(wires[716], wires[681], wires[675]);
and(wires[717], wires[682], wires[675]);
and(wires[718], wires[683], wires[675]);
and(wires[719], wires[684], wires[675]);
and(wires[720], wires[685], wires[675]);
and(wires[721], wires[686], wires[675]);
and(wires[722], wires[687], wires[675]);
not(wires[723], wires[722]);
and(wires[724], wires[680], wires[676]);
and(wires[725], wires[681], wires[676]);
and(wires[726], wires[682], wires[676]);
and(wires[727], wires[683], wires[676]);
and(wires[728], wires[684], wires[676]);
and(wires[729], wires[685], wires[676]);
and(wires[730], wires[686], wires[676]);
and(wires[731], wires[687], wires[676]);
not(wires[732], wires[731]);
and(wires[733], wires[680], wires[677]);
and(wires[734], wires[681], wires[677]);
and(wires[735], wires[682], wires[677]);
and(wires[736], wires[683], wires[677]);
and(wires[737], wires[684], wires[677]);
and(wires[738], wires[685], wires[677]);
and(wires[739], wires[686], wires[677]);
and(wires[740], wires[687], wires[677]);
not(wires[741], wires[740]);
and(wires[742], wires[680], wires[678]);
and(wires[743], wires[681], wires[678]);
and(wires[744], wires[682], wires[678]);
and(wires[745], wires[683], wires[678]);
and(wires[746], wires[684], wires[678]);
and(wires[747], wires[685], wires[678]);
and(wires[748], wires[686], wires[678]);
and(wires[749], wires[687], wires[678]);
not(wires[750], wires[749]);
and(wires[752], wires[680], wires[679]);
not(wires[753], wires[752]);
and(wires[754], wires[681], wires[679]);
not(wires[755], wires[754]);
and(wires[756], wires[682], wires[679]);
not(wires[757], wires[756]);
and(wires[758], wires[683], wires[679]);
not(wires[759], wires[758]);
and(wires[760], wires[684], wires[679]);
not(wires[761], wires[760]);
and(wires[762], wires[685], wires[679]);
not(wires[763], wires[762]);
and(wires[764], wires[686], wires[679]);
not(wires[765], wires[764]);
and(wires[766], wires[687], wires[679]);
full_adder fa_0(wires[768], wires[769], wires[16], wires[112], wires[208]);
full_adder fa_1(wires[770], wires[771], wires[304], wires[400], wires[496]);
half_adder ha_0(wires[772], wires[773], wires[592], wires[688]);
full_adder fa_2(wires[774], wires[775], wires[17], wires[25], wires[113]);
full_adder fa_3(wires[776], wires[777], wires[121], wires[209], wires[217]);
full_adder fa_4(wires[778], wires[779], wires[305], wires[313], wires[401]);
full_adder fa_5(wires[780], wires[781], wires[409], wires[497], wires[505]);
full_adder fa_6(wires[782], wires[783], wires[593], wires[601], wires[689]);
full_adder fa_7(wires[784], wires[785], wires[18], wires[26], wires[34]);
full_adder fa_8(wires[786], wires[787], wires[114], wires[122], wires[130]);
full_adder fa_9(wires[788], wires[789], wires[210], wires[218], wires[226]);
full_adder fa_10(wires[790], wires[791], wires[306], wires[314], wires[322]);
full_adder fa_11(wires[792], wires[793], wires[402], wires[410], wires[418]);
full_adder fa_12(wires[794], wires[795], wires[498], wires[506], wires[514]);
full_adder fa_13(wires[796], wires[797], wires[594], wires[602], wires[610]);
full_adder fa_14(wires[798], wires[799], wires[690], wires[698], wires[706]);
full_adder fa_15(wires[800], wires[801], wires[19], wires[27], wires[35]);
full_adder fa_16(wires[802], wires[803], wires[43], wires[115], wires[123]);
full_adder fa_17(wires[804], wires[805], wires[131], wires[139], wires[211]);
full_adder fa_18(wires[806], wires[807], wires[219], wires[227], wires[235]);
full_adder fa_19(wires[808], wires[809], wires[307], wires[315], wires[323]);
full_adder fa_20(wires[810], wires[811], wires[331], wires[403], wires[411]);
full_adder fa_21(wires[812], wires[813], wires[419], wires[427], wires[499]);
full_adder fa_22(wires[814], wires[815], wires[507], wires[515], wires[523]);
full_adder fa_23(wires[816], wires[817], wires[595], wires[603], wires[611]);
full_adder fa_24(wires[818], wires[819], wires[619], wires[691], wires[699]);
half_adder ha_1(wires[820], wires[821], wires[707], wires[715]);
full_adder fa_25(wires[822], wires[823], wires[20], wires[28], wires[36]);
full_adder fa_26(wires[824], wires[825], wires[44], wires[52], wires[116]);
full_adder fa_27(wires[826], wires[827], wires[124], wires[132], wires[140]);
full_adder fa_28(wires[828], wires[829], wires[148], wires[212], wires[220]);
full_adder fa_29(wires[830], wires[831], wires[228], wires[236], wires[244]);
full_adder fa_30(wires[832], wires[833], wires[308], wires[316], wires[324]);
full_adder fa_31(wires[834], wires[835], wires[332], wires[340], wires[404]);
full_adder fa_32(wires[836], wires[837], wires[412], wires[420], wires[428]);
full_adder fa_33(wires[838], wires[839], wires[436], wires[500], wires[508]);
full_adder fa_34(wires[840], wires[841], wires[516], wires[524], wires[532]);
full_adder fa_35(wires[842], wires[843], wires[596], wires[604], wires[612]);
full_adder fa_36(wires[844], wires[845], wires[620], wires[628], wires[692]);
full_adder fa_37(wires[846], wires[847], wires[700], wires[708], wires[716]);
full_adder fa_38(wires[848], wires[849], wires[21], wires[29], wires[37]);
full_adder fa_39(wires[850], wires[851], wires[45], wires[53], wires[61]);
full_adder fa_40(wires[852], wires[853], wires[117], wires[125], wires[133]);
full_adder fa_41(wires[854], wires[855], wires[141], wires[149], wires[157]);
full_adder fa_42(wires[856], wires[857], wires[213], wires[221], wires[229]);
full_adder fa_43(wires[858], wires[859], wires[237], wires[245], wires[253]);
full_adder fa_44(wires[860], wires[861], wires[309], wires[317], wires[325]);
full_adder fa_45(wires[862], wires[863], wires[333], wires[341], wires[349]);
full_adder fa_46(wires[864], wires[865], wires[405], wires[413], wires[421]);
full_adder fa_47(wires[866], wires[867], wires[429], wires[437], wires[445]);
full_adder fa_48(wires[868], wires[869], wires[501], wires[509], wires[517]);
full_adder fa_49(wires[870], wires[871], wires[525], wires[533], wires[541]);
full_adder fa_50(wires[872], wires[873], wires[597], wires[605], wires[613]);
full_adder fa_51(wires[874], wires[875], wires[621], wires[629], wires[637]);
full_adder fa_52(wires[876], wires[877], wires[693], wires[701], wires[709]);
full_adder fa_53(wires[878], wires[879], wires[717], wires[725], wires[733]);
full_adder fa_54(wires[880], wires[881], wires[22], wires[30], wires[38]);
full_adder fa_55(wires[882], wires[883], wires[46], wires[54], wires[62]);
full_adder fa_56(wires[884], wires[885], wires[70], wires[118], wires[126]);
full_adder fa_57(wires[886], wires[887], wires[134], wires[142], wires[150]);
full_adder fa_58(wires[888], wires[889], wires[158], wires[166], wires[214]);
full_adder fa_59(wires[890], wires[891], wires[222], wires[230], wires[238]);
full_adder fa_60(wires[892], wires[893], wires[246], wires[254], wires[262]);
full_adder fa_61(wires[894], wires[895], wires[310], wires[318], wires[326]);
full_adder fa_62(wires[896], wires[897], wires[334], wires[342], wires[350]);
full_adder fa_63(wires[898], wires[899], wires[358], wires[406], wires[414]);
full_adder fa_64(wires[900], wires[901], wires[422], wires[430], wires[438]);
full_adder fa_65(wires[902], wires[903], wires[446], wires[454], wires[502]);
full_adder fa_66(wires[904], wires[905], wires[510], wires[518], wires[526]);
full_adder fa_67(wires[906], wires[907], wires[534], wires[542], wires[550]);
full_adder fa_68(wires[908], wires[909], wires[598], wires[606], wires[614]);
full_adder fa_69(wires[910], wires[911], wires[622], wires[630], wires[638]);
full_adder fa_70(wires[912], wires[913], wires[646], wires[694], wires[702]);
full_adder fa_71(wires[914], wires[915], wires[710], wires[718], wires[726]);
half_adder ha_2(wires[916], wires[917], wires[734], wires[742]);
full_adder fa_72(wires[918], wires[919], wires[24], wires[31], wires[39]);
full_adder fa_73(wires[920], wires[921], wires[47], wires[55], wires[63]);
full_adder fa_74(wires[922], wires[923], wires[71], wires[81], wires[120]);
full_adder fa_75(wires[924], wires[925], wires[127], wires[135], wires[143]);
full_adder fa_76(wires[926], wires[927], wires[151], wires[159], wires[167]);
full_adder fa_77(wires[928], wires[929], wires[177], wires[216], wires[223]);
full_adder fa_78(wires[930], wires[931], wires[231], wires[239], wires[247]);
full_adder fa_79(wires[932], wires[933], wires[255], wires[263], wires[273]);
full_adder fa_80(wires[934], wires[935], wires[312], wires[319], wires[327]);
full_adder fa_81(wires[936], wires[937], wires[335], wires[343], wires[351]);
full_adder fa_82(wires[938], wires[939], wires[359], wires[369], wires[408]);
full_adder fa_83(wires[940], wires[941], wires[415], wires[423], wires[431]);
full_adder fa_84(wires[942], wires[943], wires[439], wires[447], wires[455]);
full_adder fa_85(wires[944], wires[945], wires[465], wires[504], wires[511]);
full_adder fa_86(wires[946], wires[947], wires[519], wires[527], wires[535]);
full_adder fa_87(wires[948], wires[949], wires[543], wires[551], wires[561]);
full_adder fa_88(wires[950], wires[951], wires[600], wires[607], wires[615]);
full_adder fa_89(wires[952], wires[953], wires[623], wires[631], wires[639]);
full_adder fa_90(wires[954], wires[955], wires[647], wires[657], wires[696]);
full_adder fa_91(wires[956], wires[957], wires[703], wires[711], wires[719]);
full_adder fa_92(wires[958], wires[959], wires[727], wires[735], wires[743]);
full_adder fa_93(wires[960], wires[961], 1'b1, wires[33], wires[40]);
full_adder fa_94(wires[962], wires[963], wires[48], wires[56], wires[64]);
full_adder fa_95(wires[964], wires[965], wires[72], wires[83], 1'b1);
full_adder fa_96(wires[966], wires[967], wires[129], wires[136], wires[144]);
full_adder fa_97(wires[968], wires[969], wires[152], wires[160], wires[168]);
full_adder fa_98(wires[970], wires[971], wires[179], 1'b1, wires[225]);
full_adder fa_99(wires[972], wires[973], wires[232], wires[240], wires[248]);
full_adder fa_100(wires[974], wires[975], wires[256], wires[264], wires[275]);
full_adder fa_101(wires[976], wires[977], 1'b1, wires[321], wires[328]);
full_adder fa_102(wires[978], wires[979], wires[336], wires[344], wires[352]);
full_adder fa_103(wires[980], wires[981], wires[360], wires[371], 1'b1);
full_adder fa_104(wires[982], wires[983], wires[417], wires[424], wires[432]);
full_adder fa_105(wires[984], wires[985], wires[440], wires[448], wires[456]);
full_adder fa_106(wires[986], wires[987], wires[467], 1'b1, wires[513]);
full_adder fa_107(wires[988], wires[989], wires[520], wires[528], wires[536]);
full_adder fa_108(wires[990], wires[991], wires[544], wires[552], wires[563]);
full_adder fa_109(wires[992], wires[993], 1'b1, wires[609], wires[616]);
full_adder fa_110(wires[994], wires[995], wires[624], wires[632], wires[640]);
full_adder fa_111(wires[996], wires[997], wires[648], wires[659], 1'b1);
full_adder fa_112(wires[998], wires[999], wires[705], wires[712], wires[720]);
full_adder fa_113(wires[1000], wires[1001], wires[728], wires[736], wires[744]);
full_adder fa_114(wires[1002], wires[1003], wires[42], wires[49], wires[57]);
full_adder fa_115(wires[1004], wires[1005], wires[65], wires[73], wires[85]);
full_adder fa_116(wires[1006], wires[1007], wires[138], wires[145], wires[153]);
full_adder fa_117(wires[1008], wires[1009], wires[161], wires[169], wires[181]);
full_adder fa_118(wires[1010], wires[1011], wires[234], wires[241], wires[249]);
full_adder fa_119(wires[1012], wires[1013], wires[257], wires[265], wires[277]);
full_adder fa_120(wires[1014], wires[1015], wires[330], wires[337], wires[345]);
full_adder fa_121(wires[1016], wires[1017], wires[353], wires[361], wires[373]);
full_adder fa_122(wires[1018], wires[1019], wires[426], wires[433], wires[441]);
full_adder fa_123(wires[1020], wires[1021], wires[449], wires[457], wires[469]);
full_adder fa_124(wires[1022], wires[1023], wires[522], wires[529], wires[537]);
full_adder fa_125(wires[1024], wires[1025], wires[545], wires[553], wires[565]);
full_adder fa_126(wires[1026], wires[1027], wires[618], wires[625], wires[633]);
full_adder fa_127(wires[1028], wires[1029], wires[641], wires[649], wires[661]);
full_adder fa_128(wires[1030], wires[1031], wires[714], wires[721], wires[729]);
full_adder fa_129(wires[1032], wires[1033], wires[737], wires[745], wires[757]);
full_adder fa_130(wires[1034], wires[1035], wires[51], wires[58], wires[66]);
full_adder fa_131(wires[1036], wires[1037], wires[74], wires[87], wires[147]);
full_adder fa_132(wires[1038], wires[1039], wires[154], wires[162], wires[170]);
full_adder fa_133(wires[1040], wires[1041], wires[183], wires[243], wires[250]);
full_adder fa_134(wires[1042], wires[1043], wires[258], wires[266], wires[279]);
full_adder fa_135(wires[1044], wires[1045], wires[339], wires[346], wires[354]);
full_adder fa_136(wires[1046], wires[1047], wires[362], wires[375], wires[435]);
full_adder fa_137(wires[1048], wires[1049], wires[442], wires[450], wires[458]);
full_adder fa_138(wires[1050], wires[1051], wires[471], wires[531], wires[538]);
full_adder fa_139(wires[1052], wires[1053], wires[546], wires[554], wires[567]);
full_adder fa_140(wires[1054], wires[1055], wires[627], wires[634], wires[642]);
full_adder fa_141(wires[1056], wires[1057], wires[650], wires[663], wires[723]);
full_adder fa_142(wires[1058], wires[1059], wires[730], wires[738], wires[746]);
full_adder fa_143(wires[1060], wires[1061], wires[60], wires[67], wires[75]);
full_adder fa_144(wires[1062], wires[1063], wires[89], wires[156], wires[163]);
full_adder fa_145(wires[1064], wires[1065], wires[171], wires[185], wires[252]);
full_adder fa_146(wires[1066], wires[1067], wires[259], wires[267], wires[281]);
full_adder fa_147(wires[1068], wires[1069], wires[348], wires[355], wires[363]);
full_adder fa_148(wires[1070], wires[1071], wires[377], wires[444], wires[451]);
full_adder fa_149(wires[1072], wires[1073], wires[459], wires[473], wires[540]);
full_adder fa_150(wires[1074], wires[1075], wires[547], wires[555], wires[569]);
full_adder fa_151(wires[1076], wires[1077], wires[636], wires[643], wires[651]);
full_adder fa_152(wires[1078], wires[1079], wires[665], wires[732], wires[739]);
half_adder ha_3(wires[1080], wires[1081], wires[747], wires[761]);
full_adder fa_153(wires[1082], wires[1083], wires[69], wires[76], wires[91]);
full_adder fa_154(wires[1084], wires[1085], wires[165], wires[172], wires[187]);
full_adder fa_155(wires[1086], wires[1087], wires[261], wires[268], wires[283]);
full_adder fa_156(wires[1088], wires[1089], wires[357], wires[364], wires[379]);
full_adder fa_157(wires[1090], wires[1091], wires[453], wires[460], wires[475]);
full_adder fa_158(wires[1092], wires[1093], wires[549], wires[556], wires[571]);
full_adder fa_159(wires[1094], wires[1095], wires[645], wires[652], wires[667]);
full_adder fa_160(wires[1096], wires[1097], wires[741], wires[748], wires[763]);
full_adder fa_161(wires[1098], wires[1099], wires[78], wires[93], wires[174]);
full_adder fa_162(wires[1100], wires[1101], wires[189], wires[270], wires[285]);
full_adder fa_163(wires[1102], wires[1103], wires[366], wires[381], wires[462]);
full_adder fa_164(wires[1104], wires[1105], wires[477], wires[558], wires[573]);
full_adder fa_165(wires[1106], wires[1107], wires[654], wires[669], wires[750]);
full_adder fa_166(wires[1108], wires[1109], wires[94], wires[190], wires[286]);
full_adder fa_167(wires[1110], wires[1111], wires[382], wires[478], wires[574]);
half_adder ha_4(wires[1112], wires[1113], wires[670], wires[766]);
full_adder fa_168(wires[1114], wires[1115], 1'b1, 1'b1, 1'b1);
full_adder fa_169(wires[1116], wires[1117], 1'b1, 1'b1, 1'b1);
half_adder ha_5(wires[1118], wires[1119], 1'b1, 1'b1);
full_adder fa_170(wires[1120], wires[1121], wires[768], wires[770], wires[772]);
full_adder fa_171(wires[1122], wires[1123], wires[769], wires[771], wires[773]);
full_adder fa_172(wires[1124], wires[1125], wires[774], wires[776], wires[778]);
full_adder fa_173(wires[1126], wires[1127], wires[780], wires[782], wires[697]);
full_adder fa_174(wires[1128], wires[1129], wires[775], wires[777], wires[779]);
full_adder fa_175(wires[1130], wires[1131], wires[781], wires[783], wires[784]);
full_adder fa_176(wires[1132], wires[1133], wires[786], wires[788], wires[790]);
full_adder fa_177(wires[1134], wires[1135], wires[792], wires[794], wires[796]);
full_adder fa_178(wires[1136], wires[1137], wires[785], wires[787], wires[789]);
full_adder fa_179(wires[1138], wires[1139], wires[791], wires[793], wires[795]);
full_adder fa_180(wires[1140], wires[1141], wires[797], wires[799], wires[800]);
full_adder fa_181(wires[1142], wires[1143], wires[802], wires[804], wires[806]);
full_adder fa_182(wires[1144], wires[1145], wires[808], wires[810], wires[812]);
full_adder fa_183(wires[1146], wires[1147], wires[814], wires[816], wires[818]);
full_adder fa_184(wires[1148], wires[1149], wires[801], wires[803], wires[805]);
full_adder fa_185(wires[1150], wires[1151], wires[807], wires[809], wires[811]);
full_adder fa_186(wires[1152], wires[1153], wires[813], wires[815], wires[817]);
full_adder fa_187(wires[1154], wires[1155], wires[819], wires[821], wires[822]);
full_adder fa_188(wires[1156], wires[1157], wires[824], wires[826], wires[828]);
full_adder fa_189(wires[1158], wires[1159], wires[830], wires[832], wires[834]);
full_adder fa_190(wires[1160], wires[1161], wires[836], wires[838], wires[840]);
full_adder fa_191(wires[1162], wires[1163], wires[842], wires[844], wires[846]);
full_adder fa_192(wires[1164], wires[1165], wires[823], wires[825], wires[827]);
full_adder fa_193(wires[1166], wires[1167], wires[829], wires[831], wires[833]);
full_adder fa_194(wires[1168], wires[1169], wires[835], wires[837], wires[839]);
full_adder fa_195(wires[1170], wires[1171], wires[841], wires[843], wires[845]);
full_adder fa_196(wires[1172], wires[1173], wires[847], wires[848], wires[850]);
full_adder fa_197(wires[1174], wires[1175], wires[852], wires[854], wires[856]);
full_adder fa_198(wires[1176], wires[1177], wires[858], wires[860], wires[862]);
full_adder fa_199(wires[1178], wires[1179], wires[864], wires[866], wires[868]);
full_adder fa_200(wires[1180], wires[1181], wires[870], wires[872], wires[874]);
half_adder ha_6(wires[1182], wires[1183], wires[876], wires[878]);
full_adder fa_201(wires[1184], wires[1185], wires[849], wires[851], wires[853]);
full_adder fa_202(wires[1186], wires[1187], wires[855], wires[857], wires[859]);
full_adder fa_203(wires[1188], wires[1189], wires[861], wires[863], wires[865]);
full_adder fa_204(wires[1190], wires[1191], wires[867], wires[869], wires[871]);
full_adder fa_205(wires[1192], wires[1193], wires[873], wires[875], wires[877]);
full_adder fa_206(wires[1194], wires[1195], wires[879], wires[880], wires[882]);
full_adder fa_207(wires[1196], wires[1197], wires[884], wires[886], wires[888]);
full_adder fa_208(wires[1198], wires[1199], wires[890], wires[892], wires[894]);
full_adder fa_209(wires[1200], wires[1201], wires[896], wires[898], wires[900]);
full_adder fa_210(wires[1202], wires[1203], wires[902], wires[904], wires[906]);
full_adder fa_211(wires[1204], wires[1205], wires[908], wires[910], wires[912]);
half_adder ha_7(wires[1206], wires[1207], wires[914], wires[916]);
full_adder fa_212(wires[1208], wires[1209], wires[881], wires[883], wires[885]);
full_adder fa_213(wires[1210], wires[1211], wires[887], wires[889], wires[891]);
full_adder fa_214(wires[1212], wires[1213], wires[893], wires[895], wires[897]);
full_adder fa_215(wires[1214], wires[1215], wires[899], wires[901], wires[903]);
full_adder fa_216(wires[1216], wires[1217], wires[905], wires[907], wires[909]);
full_adder fa_217(wires[1218], wires[1219], wires[911], wires[913], wires[915]);
full_adder fa_218(wires[1220], wires[1221], wires[917], wires[918], wires[920]);
full_adder fa_219(wires[1222], wires[1223], wires[922], wires[924], wires[926]);
full_adder fa_220(wires[1224], wires[1225], wires[928], wires[930], wires[932]);
full_adder fa_221(wires[1226], wires[1227], wires[934], wires[936], wires[938]);
full_adder fa_222(wires[1228], wires[1229], wires[940], wires[942], wires[944]);
full_adder fa_223(wires[1230], wires[1231], wires[946], wires[948], wires[950]);
full_adder fa_224(wires[1232], wires[1233], wires[952], wires[954], wires[956]);
half_adder ha_8(wires[1234], wires[1235], wires[958], wires[753]);
full_adder fa_225(wires[1236], wires[1237], wires[919], wires[921], wires[923]);
full_adder fa_226(wires[1238], wires[1239], wires[925], wires[927], wires[929]);
full_adder fa_227(wires[1240], wires[1241], wires[931], wires[933], wires[935]);
full_adder fa_228(wires[1242], wires[1243], wires[937], wires[939], wires[941]);
full_adder fa_229(wires[1244], wires[1245], wires[943], wires[945], wires[947]);
full_adder fa_230(wires[1246], wires[1247], wires[949], wires[951], wires[953]);
full_adder fa_231(wires[1248], wires[1249], wires[955], wires[957], wires[959]);
full_adder fa_232(wires[1250], wires[1251], wires[960], wires[962], wires[964]);
full_adder fa_233(wires[1252], wires[1253], wires[966], wires[968], wires[970]);
full_adder fa_234(wires[1254], wires[1255], wires[972], wires[974], wires[976]);
full_adder fa_235(wires[1256], wires[1257], wires[978], wires[980], wires[982]);
full_adder fa_236(wires[1258], wires[1259], wires[984], wires[986], wires[988]);
full_adder fa_237(wires[1260], wires[1261], wires[990], wires[992], wires[994]);
full_adder fa_238(wires[1262], wires[1263], wires[996], wires[998], wires[1000]);
full_adder fa_239(wires[1264], wires[1265], wires[961], wires[963], wires[965]);
full_adder fa_240(wires[1266], wires[1267], wires[967], wires[969], wires[971]);
full_adder fa_241(wires[1268], wires[1269], wires[973], wires[975], wires[977]);
full_adder fa_242(wires[1270], wires[1271], wires[979], wires[981], wires[983]);
full_adder fa_243(wires[1272], wires[1273], wires[985], wires[987], wires[989]);
full_adder fa_244(wires[1274], wires[1275], wires[991], wires[993], wires[995]);
full_adder fa_245(wires[1276], wires[1277], wires[997], wires[999], wires[1001]);
full_adder fa_246(wires[1278], wires[1279], wires[1002], wires[1004], wires[1006]);
full_adder fa_247(wires[1280], wires[1281], wires[1008], wires[1010], wires[1012]);
full_adder fa_248(wires[1282], wires[1283], wires[1014], wires[1016], wires[1018]);
full_adder fa_249(wires[1284], wires[1285], wires[1020], wires[1022], wires[1024]);
full_adder fa_250(wires[1286], wires[1287], wires[1026], wires[1028], wires[1030]);
full_adder fa_251(wires[1288], wires[1289], wires[1003], wires[1005], wires[1007]);
full_adder fa_252(wires[1290], wires[1291], wires[1009], wires[1011], wires[1013]);
full_adder fa_253(wires[1292], wires[1293], wires[1015], wires[1017], wires[1019]);
full_adder fa_254(wires[1294], wires[1295], wires[1021], wires[1023], wires[1025]);
full_adder fa_255(wires[1296], wires[1297], wires[1027], wires[1029], wires[1031]);
full_adder fa_256(wires[1298], wires[1299], wires[1033], wires[1034], wires[1036]);
full_adder fa_257(wires[1300], wires[1301], wires[1038], wires[1040], wires[1042]);
full_adder fa_258(wires[1302], wires[1303], wires[1044], wires[1046], wires[1048]);
full_adder fa_259(wires[1304], wires[1305], wires[1050], wires[1052], wires[1054]);
full_adder fa_260(wires[1306], wires[1307], wires[1056], wires[1058], wires[759]);
full_adder fa_261(wires[1308], wires[1309], wires[1035], wires[1037], wires[1039]);
full_adder fa_262(wires[1310], wires[1311], wires[1041], wires[1043], wires[1045]);
full_adder fa_263(wires[1312], wires[1313], wires[1047], wires[1049], wires[1051]);
full_adder fa_264(wires[1314], wires[1315], wires[1053], wires[1055], wires[1057]);
full_adder fa_265(wires[1316], wires[1317], wires[1059], wires[1060], wires[1062]);
full_adder fa_266(wires[1318], wires[1319], wires[1064], wires[1066], wires[1068]);
full_adder fa_267(wires[1320], wires[1321], wires[1070], wires[1072], wires[1074]);
full_adder fa_268(wires[1322], wires[1323], wires[1076], wires[1078], wires[1080]);
full_adder fa_269(wires[1324], wires[1325], wires[1061], wires[1063], wires[1065]);
full_adder fa_270(wires[1326], wires[1327], wires[1067], wires[1069], wires[1071]);
full_adder fa_271(wires[1328], wires[1329], wires[1073], wires[1075], wires[1077]);
full_adder fa_272(wires[1330], wires[1331], wires[1079], wires[1081], wires[1082]);
full_adder fa_273(wires[1332], wires[1333], wires[1084], wires[1086], wires[1088]);
full_adder fa_274(wires[1334], wires[1335], wires[1090], wires[1092], wires[1094]);
full_adder fa_275(wires[1336], wires[1337], wires[1083], wires[1085], wires[1087]);
full_adder fa_276(wires[1338], wires[1339], wires[1089], wires[1091], wires[1093]);
full_adder fa_277(wires[1340], wires[1341], wires[1095], wires[1097], wires[1098]);
full_adder fa_278(wires[1342], wires[1343], wires[1100], wires[1102], wires[1104]);
half_adder ha_9(wires[1344], wires[1345], wires[1106], wires[765]);
full_adder fa_279(wires[1346], wires[1347], wires[1099], wires[1101], wires[1103]);
full_adder fa_280(wires[1348], wires[1349], wires[1105], wires[1107], wires[1108]);
half_adder ha_10(wires[1350], wires[1351], wires[1110], wires[1112]);
full_adder fa_281(wires[1352], wires[1353], wires[1109], wires[1111], wires[1113]);
full_adder fa_282(wires[1354], wires[1355], wires[1114], wires[1116], wires[1118]);
full_adder fa_283(wires[1356], wires[1357], wires[1115], wires[1117], wires[1119]);
full_adder fa_284(wires[1358], wires[1359], wires[1121], wires[1122], wires[1124]);
full_adder fa_285(wires[1360], wires[1361], wires[1123], wires[1125], wires[1127]);
full_adder fa_286(wires[1362], wires[1363], wires[1128], wires[1130], wires[1132]);
half_adder ha_11(wires[1364], wires[1365], wires[1134], wires[798]);
full_adder fa_287(wires[1366], wires[1367], wires[1129], wires[1131], wires[1133]);
full_adder fa_288(wires[1368], wires[1369], wires[1135], wires[1136], wires[1138]);
full_adder fa_289(wires[1370], wires[1371], wires[1140], wires[1142], wires[1144]);
half_adder ha_12(wires[1372], wires[1373], wires[1146], wires[820]);
full_adder fa_290(wires[1374], wires[1375], wires[1137], wires[1139], wires[1141]);
full_adder fa_291(wires[1376], wires[1377], wires[1143], wires[1145], wires[1147]);
full_adder fa_292(wires[1378], wires[1379], wires[1148], wires[1150], wires[1152]);
full_adder fa_293(wires[1380], wires[1381], wires[1154], wires[1156], wires[1158]);
full_adder fa_294(wires[1382], wires[1383], wires[1160], wires[1162], wires[724]);
full_adder fa_295(wires[1384], wires[1385], wires[1149], wires[1151], wires[1153]);
full_adder fa_296(wires[1386], wires[1387], wires[1155], wires[1157], wires[1159]);
full_adder fa_297(wires[1388], wires[1389], wires[1161], wires[1163], wires[1164]);
full_adder fa_298(wires[1390], wires[1391], wires[1166], wires[1168], wires[1170]);
full_adder fa_299(wires[1392], wires[1393], wires[1172], wires[1174], wires[1176]);
full_adder fa_300(wires[1394], wires[1395], wires[1178], wires[1180], wires[1182]);
full_adder fa_301(wires[1396], wires[1397], wires[1165], wires[1167], wires[1169]);
full_adder fa_302(wires[1398], wires[1399], wires[1171], wires[1173], wires[1175]);
full_adder fa_303(wires[1400], wires[1401], wires[1177], wires[1179], wires[1181]);
full_adder fa_304(wires[1402], wires[1403], wires[1183], wires[1184], wires[1186]);
full_adder fa_305(wires[1404], wires[1405], wires[1188], wires[1190], wires[1192]);
full_adder fa_306(wires[1406], wires[1407], wires[1194], wires[1196], wires[1198]);
full_adder fa_307(wires[1408], wires[1409], wires[1200], wires[1202], wires[1204]);
full_adder fa_308(wires[1410], wires[1411], wires[1185], wires[1187], wires[1189]);
full_adder fa_309(wires[1412], wires[1413], wires[1191], wires[1193], wires[1195]);
full_adder fa_310(wires[1414], wires[1415], wires[1197], wires[1199], wires[1201]);
full_adder fa_311(wires[1416], wires[1417], wires[1203], wires[1205], wires[1207]);
full_adder fa_312(wires[1418], wires[1419], wires[1208], wires[1210], wires[1212]);
full_adder fa_313(wires[1420], wires[1421], wires[1214], wires[1216], wires[1218]);
full_adder fa_314(wires[1422], wires[1423], wires[1220], wires[1222], wires[1224]);
full_adder fa_315(wires[1424], wires[1425], wires[1226], wires[1228], wires[1230]);
half_adder ha_13(wires[1426], wires[1427], wires[1232], wires[1234]);
full_adder fa_316(wires[1428], wires[1429], wires[1209], wires[1211], wires[1213]);
full_adder fa_317(wires[1430], wires[1431], wires[1215], wires[1217], wires[1219]);
full_adder fa_318(wires[1432], wires[1433], wires[1221], wires[1223], wires[1225]);
full_adder fa_319(wires[1434], wires[1435], wires[1227], wires[1229], wires[1231]);
full_adder fa_320(wires[1436], wires[1437], wires[1233], wires[1235], wires[1236]);
full_adder fa_321(wires[1438], wires[1439], wires[1238], wires[1240], wires[1242]);
full_adder fa_322(wires[1440], wires[1441], wires[1244], wires[1246], wires[1248]);
full_adder fa_323(wires[1442], wires[1443], wires[1250], wires[1252], wires[1254]);
full_adder fa_324(wires[1444], wires[1445], wires[1256], wires[1258], wires[1260]);
half_adder ha_14(wires[1446], wires[1447], wires[1262], wires[755]);
full_adder fa_325(wires[1448], wires[1449], wires[1237], wires[1239], wires[1241]);
full_adder fa_326(wires[1450], wires[1451], wires[1243], wires[1245], wires[1247]);
full_adder fa_327(wires[1452], wires[1453], wires[1249], wires[1251], wires[1253]);
full_adder fa_328(wires[1454], wires[1455], wires[1255], wires[1257], wires[1259]);
full_adder fa_329(wires[1456], wires[1457], wires[1261], wires[1263], wires[1264]);
full_adder fa_330(wires[1458], wires[1459], wires[1266], wires[1268], wires[1270]);
full_adder fa_331(wires[1460], wires[1461], wires[1272], wires[1274], wires[1276]);
full_adder fa_332(wires[1462], wires[1463], wires[1278], wires[1280], wires[1282]);
full_adder fa_333(wires[1464], wires[1465], wires[1284], wires[1286], wires[1032]);
full_adder fa_334(wires[1466], wires[1467], wires[1265], wires[1267], wires[1269]);
full_adder fa_335(wires[1468], wires[1469], wires[1271], wires[1273], wires[1275]);
full_adder fa_336(wires[1470], wires[1471], wires[1277], wires[1279], wires[1281]);
full_adder fa_337(wires[1472], wires[1473], wires[1283], wires[1285], wires[1287]);
full_adder fa_338(wires[1474], wires[1475], wires[1288], wires[1290], wires[1292]);
full_adder fa_339(wires[1476], wires[1477], wires[1294], wires[1296], wires[1298]);
full_adder fa_340(wires[1478], wires[1479], wires[1300], wires[1302], wires[1304]);
full_adder fa_341(wires[1480], wires[1481], wires[1289], wires[1291], wires[1293]);
full_adder fa_342(wires[1482], wires[1483], wires[1295], wires[1297], wires[1299]);
full_adder fa_343(wires[1484], wires[1485], wires[1301], wires[1303], wires[1305]);
full_adder fa_344(wires[1486], wires[1487], wires[1307], wires[1308], wires[1310]);
full_adder fa_345(wires[1488], wires[1489], wires[1312], wires[1314], wires[1316]);
full_adder fa_346(wires[1490], wires[1491], wires[1318], wires[1320], wires[1322]);
full_adder fa_347(wires[1492], wires[1493], wires[1309], wires[1311], wires[1313]);
full_adder fa_348(wires[1494], wires[1495], wires[1315], wires[1317], wires[1319]);
full_adder fa_349(wires[1496], wires[1497], wires[1321], wires[1323], wires[1324]);
full_adder fa_350(wires[1498], wires[1499], wires[1326], wires[1328], wires[1330]);
full_adder fa_351(wires[1500], wires[1501], wires[1332], wires[1334], wires[1096]);
full_adder fa_352(wires[1502], wires[1503], wires[1325], wires[1327], wires[1329]);
full_adder fa_353(wires[1504], wires[1505], wires[1331], wires[1333], wires[1335]);
full_adder fa_354(wires[1506], wires[1507], wires[1336], wires[1338], wires[1340]);
half_adder ha_15(wires[1508], wires[1509], wires[1342], wires[1344]);
full_adder fa_355(wires[1510], wires[1511], wires[1337], wires[1339], wires[1341]);
full_adder fa_356(wires[1512], wires[1513], wires[1343], wires[1345], wires[1346]);
half_adder ha_16(wires[1514], wires[1515], wires[1348], wires[1350]);
full_adder fa_357(wires[1516], wires[1517], wires[1347], wires[1349], wires[1351]);
half_adder ha_17(wires[1518], wires[1519], wires[1352], wires[1354]);
full_adder fa_358(wires[1520], wires[1521], wires[1353], wires[1355], wires[1356]);
half_adder ha_18(wires[1522], wires[1523], wires[1358], wires[1126]);
full_adder fa_359(wires[1524], wires[1525], wires[1359], wires[1360], wires[1362]);
full_adder fa_360(wires[1526], wires[1527], wires[1361], wires[1363], wires[1365]);
full_adder fa_361(wires[1528], wires[1529], wires[1366], wires[1368], wires[1370]);
full_adder fa_362(wires[1530], wires[1531], wires[1367], wires[1369], wires[1371]);
full_adder fa_363(wires[1532], wires[1533], wires[1373], wires[1374], wires[1376]);
full_adder fa_364(wires[1534], wires[1535], wires[1378], wires[1380], wires[1382]);
full_adder fa_365(wires[1536], wires[1537], wires[1375], wires[1377], wires[1379]);
full_adder fa_366(wires[1538], wires[1539], wires[1381], wires[1383], wires[1384]);
full_adder fa_367(wires[1540], wires[1541], wires[1386], wires[1388], wires[1390]);
half_adder ha_19(wires[1542], wires[1543], wires[1392], wires[1394]);
full_adder fa_368(wires[1544], wires[1545], wires[1385], wires[1387], wires[1389]);
full_adder fa_369(wires[1546], wires[1547], wires[1391], wires[1393], wires[1395]);
full_adder fa_370(wires[1548], wires[1549], wires[1396], wires[1398], wires[1400]);
full_adder fa_371(wires[1550], wires[1551], wires[1402], wires[1404], wires[1406]);
half_adder ha_20(wires[1552], wires[1553], wires[1408], wires[1206]);
full_adder fa_372(wires[1554], wires[1555], wires[1397], wires[1399], wires[1401]);
full_adder fa_373(wires[1556], wires[1557], wires[1403], wires[1405], wires[1407]);
full_adder fa_374(wires[1558], wires[1559], wires[1409], wires[1410], wires[1412]);
full_adder fa_375(wires[1560], wires[1561], wires[1414], wires[1416], wires[1418]);
full_adder fa_376(wires[1562], wires[1563], wires[1420], wires[1422], wires[1424]);
full_adder fa_377(wires[1564], wires[1565], wires[1411], wires[1413], wires[1415]);
full_adder fa_378(wires[1566], wires[1567], wires[1417], wires[1419], wires[1421]);
full_adder fa_379(wires[1568], wires[1569], wires[1423], wires[1425], wires[1427]);
full_adder fa_380(wires[1570], wires[1571], wires[1428], wires[1430], wires[1432]);
full_adder fa_381(wires[1572], wires[1573], wires[1434], wires[1436], wires[1438]);
full_adder fa_382(wires[1574], wires[1575], wires[1440], wires[1442], wires[1444]);
full_adder fa_383(wires[1576], wires[1577], wires[1429], wires[1431], wires[1433]);
full_adder fa_384(wires[1578], wires[1579], wires[1435], wires[1437], wires[1439]);
full_adder fa_385(wires[1580], wires[1581], wires[1441], wires[1443], wires[1445]);
full_adder fa_386(wires[1582], wires[1583], wires[1447], wires[1448], wires[1450]);
full_adder fa_387(wires[1584], wires[1585], wires[1452], wires[1454], wires[1456]);
full_adder fa_388(wires[1586], wires[1587], wires[1458], wires[1460], wires[1462]);
full_adder fa_389(wires[1588], wires[1589], wires[1449], wires[1451], wires[1453]);
full_adder fa_390(wires[1590], wires[1591], wires[1455], wires[1457], wires[1459]);
full_adder fa_391(wires[1592], wires[1593], wires[1461], wires[1463], wires[1465]);
full_adder fa_392(wires[1594], wires[1595], wires[1466], wires[1468], wires[1470]);
full_adder fa_393(wires[1596], wires[1597], wires[1472], wires[1474], wires[1476]);
half_adder ha_21(wires[1598], wires[1599], wires[1478], wires[1306]);
full_adder fa_394(wires[1600], wires[1601], wires[1467], wires[1469], wires[1471]);
full_adder fa_395(wires[1602], wires[1603], wires[1473], wires[1475], wires[1477]);
full_adder fa_396(wires[1604], wires[1605], wires[1479], wires[1480], wires[1482]);
full_adder fa_397(wires[1606], wires[1607], wires[1484], wires[1486], wires[1488]);
full_adder fa_398(wires[1608], wires[1609], wires[1481], wires[1483], wires[1485]);
full_adder fa_399(wires[1610], wires[1611], wires[1487], wires[1489], wires[1491]);
full_adder fa_400(wires[1612], wires[1613], wires[1492], wires[1494], wires[1496]);
half_adder ha_22(wires[1614], wires[1615], wires[1498], wires[1500]);
full_adder fa_401(wires[1616], wires[1617], wires[1493], wires[1495], wires[1497]);
full_adder fa_402(wires[1618], wires[1619], wires[1499], wires[1501], wires[1502]);
full_adder fa_403(wires[1620], wires[1621], wires[1504], wires[1506], wires[1508]);
full_adder fa_404(wires[1622], wires[1623], wires[1503], wires[1505], wires[1507]);
full_adder fa_405(wires[1624], wires[1625], wires[1509], wires[1510], wires[1512]);
full_adder fa_406(wires[1626], wires[1627], wires[1511], wires[1513], wires[1515]);
half_adder ha_23(wires[1628], wires[1629], wires[1516], wires[1518]);
full_adder fa_407(wires[1630], wires[1631], wires[1517], wires[1519], wires[1520]);
half_adder ha_24(wires[1632], wires[1633], wires[1521], wires[1357]);
full_adder fa_408(wires[1634], wires[1635], wires[1523], wires[1524], wires[1364]);
full_adder fa_409(wires[1636], wires[1637], wires[1525], wires[1526], wires[1528]);
full_adder fa_410(wires[1638], wires[1639], wires[1527], wires[1529], wires[1530]);
half_adder ha_25(wires[1640], wires[1641], wires[1532], wires[1534]);
full_adder fa_411(wires[1642], wires[1643], wires[1531], wires[1533], wires[1535]);
full_adder fa_412(wires[1644], wires[1645], wires[1536], wires[1538], wires[1540]);
full_adder fa_413(wires[1646], wires[1647], wires[1537], wires[1539], wires[1541]);
full_adder fa_414(wires[1648], wires[1649], wires[1543], wires[1544], wires[1546]);
full_adder fa_415(wires[1650], wires[1651], wires[1548], wires[1550], wires[1552]);
full_adder fa_416(wires[1652], wires[1653], wires[1545], wires[1547], wires[1549]);
full_adder fa_417(wires[1654], wires[1655], wires[1551], wires[1553], wires[1554]);
full_adder fa_418(wires[1656], wires[1657], wires[1556], wires[1558], wires[1560]);
half_adder ha_26(wires[1658], wires[1659], wires[1562], wires[1426]);
full_adder fa_419(wires[1660], wires[1661], wires[1555], wires[1557], wires[1559]);
full_adder fa_420(wires[1662], wires[1663], wires[1561], wires[1563], wires[1564]);
full_adder fa_421(wires[1664], wires[1665], wires[1566], wires[1568], wires[1570]);
full_adder fa_422(wires[1666], wires[1667], wires[1572], wires[1574], wires[1446]);
full_adder fa_423(wires[1668], wires[1669], wires[1565], wires[1567], wires[1569]);
full_adder fa_424(wires[1670], wires[1671], wires[1571], wires[1573], wires[1575]);
full_adder fa_425(wires[1672], wires[1673], wires[1576], wires[1578], wires[1580]);
full_adder fa_426(wires[1674], wires[1675], wires[1582], wires[1584], wires[1586]);
full_adder fa_427(wires[1676], wires[1677], wires[1577], wires[1579], wires[1581]);
full_adder fa_428(wires[1678], wires[1679], wires[1583], wires[1585], wires[1587]);
full_adder fa_429(wires[1680], wires[1681], wires[1588], wires[1590], wires[1592]);
full_adder fa_430(wires[1682], wires[1683], wires[1594], wires[1596], wires[1598]);
full_adder fa_431(wires[1684], wires[1685], wires[1589], wires[1591], wires[1593]);
full_adder fa_432(wires[1686], wires[1687], wires[1595], wires[1597], wires[1599]);
full_adder fa_433(wires[1688], wires[1689], wires[1600], wires[1602], wires[1604]);
half_adder ha_27(wires[1690], wires[1691], wires[1606], wires[1490]);
full_adder fa_434(wires[1692], wires[1693], wires[1601], wires[1603], wires[1605]);
full_adder fa_435(wires[1694], wires[1695], wires[1607], wires[1608], wires[1610]);
half_adder ha_28(wires[1696], wires[1697], wires[1612], wires[1614]);
full_adder fa_436(wires[1698], wires[1699], wires[1609], wires[1611], wires[1613]);
full_adder fa_437(wires[1700], wires[1701], wires[1615], wires[1616], wires[1618]);
full_adder fa_438(wires[1702], wires[1703], wires[1617], wires[1619], wires[1621]);
full_adder fa_439(wires[1704], wires[1705], wires[1622], wires[1624], wires[1514]);
full_adder fa_440(wires[1706], wires[1707], wires[1623], wires[1625], wires[1626]);
full_adder fa_441(wires[1708], wires[1709], wires[1627], wires[1629], wires[1630]);
half_adder ha_29(wires[1710], wires[1711], wires[1631], wires[1632]);
full_adder fa_442(wires[1712], wires[1713], wires[1635], wires[1636], wires[1372]);
full_adder fa_443(wires[1714], wires[1715], wires[1637], wires[1638], wires[1640]);
full_adder fa_444(wires[1716], wires[1717], wires[1639], wires[1641], wires[1642]);
half_adder ha_30(wires[1718], wires[1719], wires[1644], wires[1542]);
full_adder fa_445(wires[1720], wires[1721], wires[1643], wires[1645], wires[1646]);
half_adder ha_31(wires[1722], wires[1723], wires[1648], wires[1650]);
full_adder fa_446(wires[1724], wires[1725], wires[1647], wires[1649], wires[1651]);
full_adder fa_447(wires[1726], wires[1727], wires[1652], wires[1654], wires[1656]);
full_adder fa_448(wires[1728], wires[1729], wires[1653], wires[1655], wires[1657]);
full_adder fa_449(wires[1730], wires[1731], wires[1659], wires[1660], wires[1662]);
half_adder ha_32(wires[1732], wires[1733], wires[1664], wires[1666]);
full_adder fa_450(wires[1734], wires[1735], wires[1661], wires[1663], wires[1665]);
full_adder fa_451(wires[1736], wires[1737], wires[1667], wires[1668], wires[1670]);
full_adder fa_452(wires[1738], wires[1739], wires[1672], wires[1674], wires[1464]);
full_adder fa_453(wires[1740], wires[1741], wires[1669], wires[1671], wires[1673]);
full_adder fa_454(wires[1742], wires[1743], wires[1675], wires[1676], wires[1678]);
half_adder ha_33(wires[1744], wires[1745], wires[1680], wires[1682]);
full_adder fa_455(wires[1746], wires[1747], wires[1677], wires[1679], wires[1681]);
full_adder fa_456(wires[1748], wires[1749], wires[1683], wires[1684], wires[1686]);
half_adder ha_34(wires[1750], wires[1751], wires[1688], wires[1690]);
full_adder fa_457(wires[1752], wires[1753], wires[1685], wires[1687], wires[1689]);
full_adder fa_458(wires[1754], wires[1755], wires[1691], wires[1692], wires[1694]);
full_adder fa_459(wires[1756], wires[1757], wires[1693], wires[1695], wires[1697]);
full_adder fa_460(wires[1758], wires[1759], wires[1698], wires[1700], wires[1620]);
full_adder fa_461(wires[1760], wires[1761], wires[1699], wires[1701], wires[1702]);
full_adder fa_462(wires[1762], wires[1763], wires[1703], wires[1705], wires[1706]);
half_adder ha_35(wires[1764], wires[1765], wires[1707], wires[1708]);
half_adder ha_36(wires[1766], wires[1767], wires[1709], wires[1710]);
half_adder ha_37(wires[1768], wires[1769], wires[1711], wires[1633]);
half_adder ha_38(wires[1770], wires[1771], wires[1713], wires[1714]);
full_adder fa_463(wires[1772], wires[1773], wires[1715], wires[1716], wires[1718]);
full_adder fa_464(wires[1774], wires[1775], wires[1717], wires[1719], wires[1720]);
full_adder fa_465(wires[1776], wires[1777], wires[1721], wires[1723], wires[1724]);
half_adder ha_39(wires[1778], wires[1779], wires[1726], wires[1658]);
full_adder fa_466(wires[1780], wires[1781], wires[1725], wires[1727], wires[1728]);
half_adder ha_40(wires[1782], wires[1783], wires[1730], wires[1732]);
full_adder fa_467(wires[1784], wires[1785], wires[1729], wires[1731], wires[1733]);
full_adder fa_468(wires[1786], wires[1787], wires[1734], wires[1736], wires[1738]);
full_adder fa_469(wires[1788], wires[1789], wires[1735], wires[1737], wires[1739]);
full_adder fa_470(wires[1790], wires[1791], wires[1740], wires[1742], wires[1744]);
full_adder fa_471(wires[1792], wires[1793], wires[1741], wires[1743], wires[1745]);
full_adder fa_472(wires[1794], wires[1795], wires[1746], wires[1748], wires[1750]);
full_adder fa_473(wires[1796], wires[1797], wires[1747], wires[1749], wires[1751]);
full_adder fa_474(wires[1798], wires[1799], wires[1752], wires[1754], wires[1696]);
full_adder fa_475(wires[1800], wires[1801], wires[1753], wires[1755], wires[1756]);
full_adder fa_476(wires[1802], wires[1803], wires[1757], wires[1759], wires[1760]);
full_adder fa_477(wires[1804], wires[1805], wires[1761], wires[1762], wires[1628]);
half_adder ha_41(wires[1806], wires[1807], wires[1763], wires[1764]);
half_adder ha_42(wires[1808], wires[1809], wires[1765], wires[1766]);
half_adder ha_43(wires[1810], wires[1811], wires[1767], wires[1768]);
half_adder ha_44(wires[1812], wires[1813], wires[1771], wires[1772]);
full_adder fa_478(wires[1814], wires[1815], wires[1773], wires[1774], wires[1722]);
full_adder fa_479(wires[1816], wires[1817], wires[1775], wires[1776], wires[1778]);
full_adder fa_480(wires[1818], wires[1819], wires[1777], wires[1779], wires[1780]);
full_adder fa_481(wires[1820], wires[1821], wires[1781], wires[1783], wires[1784]);
full_adder fa_482(wires[1822], wires[1823], wires[1785], wires[1787], wires[1788]);
full_adder fa_483(wires[1824], wires[1825], wires[1789], wires[1791], wires[1792]);
full_adder fa_484(wires[1826], wires[1827], wires[1793], wires[1795], wires[1796]);
full_adder fa_485(wires[1828], wires[1829], wires[1797], wires[1799], wires[1800]);
full_adder fa_486(wires[1830], wires[1831], wires[1801], wires[1802], wires[1704]);
half_adder ha_45(wires[1832], wires[1833], wires[1803], wires[1804]);
half_adder ha_46(wires[1834], wires[1835], wires[1805], wires[1806]);
half_adder ha_47(wires[1836], wires[1837], wires[1807], wires[1808]);
half_adder ha_48(wires[1838], wires[1839], wires[1809], wires[1810]);
half_adder ha_49(wires[1840], wires[1841], wires[1811], wires[1769]);
half_adder ha_50(wires[1842], wires[1843], wires[1813], wires[1814]);
half_adder ha_51(wires[1844], wires[1845], wires[1815], wires[1816]);
full_adder fa_487(wires[1846], wires[1847], wires[1817], wires[1818], wires[1782]);
full_adder fa_488(wires[1848], wires[1849], wires[1819], wires[1820], wires[1786]);
full_adder fa_489(wires[1850], wires[1851], wires[1821], wires[1822], wires[1790]);
full_adder fa_490(wires[1852], wires[1853], wires[1823], wires[1824], wires[1794]);
full_adder fa_491(wires[1854], wires[1855], wires[1825], wires[1826], wires[1798]);
full_adder fa_492(wires[1856], wires[1857], wires[1827], wires[1828], wires[1758]);
half_adder ha_52(wires[1858], wires[1859], wires[1829], wires[1830]);
half_adder ha_53(wires[1860], wires[1861], wires[1831], wires[1832]);
half_adder ha_54(wires[1862], wires[1863], wires[1833], wires[1834]);
half_adder ha_55(wires[1864], wires[1865], wires[1835], wires[1836]);
half_adder ha_56(wires[1866], wires[1867], wires[1837], wires[1838]);
half_adder ha_57(wires[1868], wires[1869], wires[1839], wires[1840]);
half_adder ha_58(wires[1870], wires[1871], wires[1843], wires[1844]);
full_adder fa_493(wires[1872], wires[1873], wires[1845], wires[1846], wires[1871]);
full_adder fa_494(wires[1874], wires[1875], wires[1847], wires[1848], wires[1873]);
full_adder fa_495(wires[1876], wires[1877], wires[1849], wires[1850], wires[1875]);
full_adder fa_496(wires[1878], wires[1879], wires[1851], wires[1852], wires[1877]);
full_adder fa_497(wires[1880], wires[1881], wires[1853], wires[1854], wires[1879]);
full_adder fa_498(wires[1882], wires[1883], wires[1855], wires[1856], wires[1881]);
full_adder fa_499(wires[1884], wires[1885], wires[1857], wires[1858], wires[1883]);
full_adder fa_500(wires[1886], wires[1887], wires[1859], wires[1860], wires[1885]);
full_adder fa_501(wires[1888], wires[1889], wires[1861], wires[1862], wires[1887]);
full_adder fa_502(wires[1890], wires[1891], wires[1863], wires[1864], wires[1889]);
full_adder fa_503(wires[1892], wires[1893], wires[1865], wires[1866], wires[1891]);
full_adder fa_504(wires[1894], wires[1895], wires[1867], wires[1868], wires[1893]);
full_adder fa_505(wires[1896], wires[1897], wires[1869], wires[1841], wires[1895]);
endmodule