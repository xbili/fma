module fma_4x4(out_0, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7);
input [3:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
output [9:0] out_0;
wire [257:0] wires;
assign wires[0] = in_0[0];
assign wires[1] = in_0[1];
assign wires[2] = in_0[2];
assign wires[3] = in_0[3];
assign wires[4] = in_1[0];
assign wires[5] = in_1[1];
assign wires[6] = in_1[2];
assign wires[7] = in_1[3];
assign wires[30] = in_2[0];
assign wires[31] = in_2[1];
assign wires[32] = in_2[2];
assign wires[33] = in_2[3];
assign wires[34] = in_3[0];
assign wires[35] = in_3[1];
assign wires[36] = in_3[2];
assign wires[37] = in_3[3];
assign wires[60] = in_4[0];
assign wires[61] = in_4[1];
assign wires[62] = in_4[2];
assign wires[63] = in_4[3];
assign wires[64] = in_5[0];
assign wires[65] = in_5[1];
assign wires[66] = in_5[2];
assign wires[67] = in_5[3];
assign wires[90] = in_6[0];
assign wires[91] = in_6[1];
assign wires[92] = in_6[2];
assign wires[93] = in_6[3];
assign wires[94] = in_7[0];
assign wires[95] = in_7[1];
assign wires[96] = in_7[2];
assign wires[97] = in_7[3];
assign out_0[0] = wires[166];
assign out_0[1] = wires[196];
assign out_0[2] = wires[216];
assign out_0[3] = wires[230];
assign out_0[4] = wires[244];
assign out_0[5] = wires[246];
assign out_0[6] = wires[248];
assign out_0[7] = wires[250];
assign out_0[8] = wires[252];
assign out_0[9] = wires[254];
and(wires[8], wires[4], wires[0]);
and(wires[9], wires[5], wires[0]);
and(wires[10], wires[6], wires[0]);
and(wires[11], wires[7], wires[0]);
not(wires[12], wires[11]);
and(wires[13], wires[4], wires[1]);
and(wires[14], wires[5], wires[1]);
and(wires[15], wires[6], wires[1]);
and(wires[16], wires[7], wires[1]);
not(wires[17], wires[16]);
and(wires[18], wires[4], wires[2]);
and(wires[19], wires[5], wires[2]);
and(wires[20], wires[6], wires[2]);
and(wires[21], wires[7], wires[2]);
not(wires[22], wires[21]);
and(wires[23], wires[4], wires[3]);
not(wires[24], wires[23]);
and(wires[25], wires[5], wires[3]);
not(wires[26], wires[25]);
and(wires[27], wires[6], wires[3]);
not(wires[28], wires[27]);
and(wires[29], wires[7], wires[3]);
and(wires[38], wires[34], wires[30]);
and(wires[39], wires[35], wires[30]);
and(wires[40], wires[36], wires[30]);
and(wires[41], wires[37], wires[30]);
not(wires[42], wires[41]);
and(wires[43], wires[34], wires[31]);
and(wires[44], wires[35], wires[31]);
and(wires[45], wires[36], wires[31]);
and(wires[46], wires[37], wires[31]);
not(wires[47], wires[46]);
and(wires[48], wires[34], wires[32]);
and(wires[49], wires[35], wires[32]);
and(wires[50], wires[36], wires[32]);
and(wires[51], wires[37], wires[32]);
not(wires[52], wires[51]);
and(wires[53], wires[34], wires[33]);
not(wires[54], wires[53]);
and(wires[55], wires[35], wires[33]);
not(wires[56], wires[55]);
and(wires[57], wires[36], wires[33]);
not(wires[58], wires[57]);
and(wires[59], wires[37], wires[33]);
and(wires[68], wires[64], wires[60]);
and(wires[69], wires[65], wires[60]);
and(wires[70], wires[66], wires[60]);
and(wires[71], wires[67], wires[60]);
not(wires[72], wires[71]);
and(wires[73], wires[64], wires[61]);
and(wires[74], wires[65], wires[61]);
and(wires[75], wires[66], wires[61]);
and(wires[76], wires[67], wires[61]);
not(wires[77], wires[76]);
and(wires[78], wires[64], wires[62]);
and(wires[79], wires[65], wires[62]);
and(wires[80], wires[66], wires[62]);
and(wires[81], wires[67], wires[62]);
not(wires[82], wires[81]);
and(wires[83], wires[64], wires[63]);
not(wires[84], wires[83]);
and(wires[85], wires[65], wires[63]);
not(wires[86], wires[85]);
and(wires[87], wires[66], wires[63]);
not(wires[88], wires[87]);
and(wires[89], wires[67], wires[63]);
and(wires[98], wires[94], wires[90]);
and(wires[99], wires[95], wires[90]);
and(wires[100], wires[96], wires[90]);
and(wires[101], wires[97], wires[90]);
not(wires[102], wires[101]);
and(wires[103], wires[94], wires[91]);
and(wires[104], wires[95], wires[91]);
and(wires[105], wires[96], wires[91]);
and(wires[106], wires[97], wires[91]);
not(wires[107], wires[106]);
and(wires[108], wires[94], wires[92]);
and(wires[109], wires[95], wires[92]);
and(wires[110], wires[96], wires[92]);
and(wires[111], wires[97], wires[92]);
not(wires[112], wires[111]);
and(wires[113], wires[94], wires[93]);
not(wires[114], wires[113]);
and(wires[115], wires[95], wires[93]);
not(wires[116], wires[115]);
and(wires[117], wires[96], wires[93]);
not(wires[118], wires[117]);
and(wires[119], wires[97], wires[93]);
full_adder fa_0(wires[122], wires[123], wires[8], wires[38], wires[68]);
full_adder fa_1(wires[124], wires[125], wires[9], wires[13], wires[39]);
full_adder fa_2(wires[126], wires[127], wires[43], wires[69], wires[73]);
half_adder ha_0(wires[128], wires[129], wires[99], wires[103]);
full_adder fa_3(wires[130], wires[131], wires[10], wires[14], wires[18]);
full_adder fa_4(wires[132], wires[133], wires[40], wires[44], wires[48]);
full_adder fa_5(wires[134], wires[135], wires[70], wires[74], wires[78]);
full_adder fa_6(wires[136], wires[137], wires[100], wires[104], wires[108]);
full_adder fa_7(wires[138], wires[139], wires[12], wires[15], wires[19]);
full_adder fa_8(wires[140], wires[141], wires[24], wires[42], wires[45]);
full_adder fa_9(wires[142], wires[143], wires[49], wires[54], wires[72]);
full_adder fa_10(wires[144], wires[145], wires[75], wires[79], wires[84]);
full_adder fa_11(wires[146], wires[147], wires[102], wires[105], wires[109]);
full_adder fa_12(wires[148], wires[149], wires[17], wires[20], wires[26]);
full_adder fa_13(wires[150], wires[151], wires[47], wires[50], wires[56]);
full_adder fa_14(wires[152], wires[153], wires[77], wires[80], wires[86]);
full_adder fa_15(wires[154], wires[155], wires[107], wires[110], wires[116]);
full_adder fa_16(wires[156], wires[157], wires[22], wires[28], wires[52]);
full_adder fa_17(wires[158], wires[159], wires[58], wires[82], wires[88]);
half_adder ha_1(wires[160], wires[161], wires[112], wires[118]);
full_adder fa_18(wires[162], wires[163], wires[29], wires[59], wires[89]);
half_adder ha_2(wires[164], wires[165], wires[119], 1'b1);
half_adder ha_3(wires[166], wires[167], wires[122], wires[98]);
full_adder fa_19(wires[168], wires[169], wires[123], wires[124], wires[126]);
full_adder fa_20(wires[170], wires[171], wires[125], wires[127], wires[129]);
full_adder fa_21(wires[172], wires[173], wires[130], wires[132], wires[134]);
full_adder fa_22(wires[174], wires[175], wires[131], wires[133], wires[135]);
full_adder fa_23(wires[176], wires[177], wires[137], wires[138], wires[140]);
full_adder fa_24(wires[178], wires[179], wires[142], wires[144], wires[146]);
full_adder fa_25(wires[180], wires[181], wires[139], wires[141], wires[143]);
full_adder fa_26(wires[182], wires[183], wires[145], wires[147], wires[148]);
full_adder fa_27(wires[184], wires[185], wires[150], wires[152], wires[154]);
full_adder fa_28(wires[186], wires[187], wires[149], wires[151], wires[153]);
full_adder fa_29(wires[188], wires[189], wires[155], wires[156], wires[158]);
full_adder fa_30(wires[190], wires[191], wires[157], wires[159], wires[161]);
half_adder ha_4(wires[192], wires[193], wires[162], wires[164]);
half_adder ha_5(wires[194], wires[195], wires[163], wires[165]);
full_adder fa_31(wires[196], wires[197], wires[167], wires[168], wires[128]);
full_adder fa_32(wires[198], wires[199], wires[169], wires[170], wires[172]);
full_adder fa_33(wires[200], wires[201], wires[171], wires[173], wires[174]);
full_adder fa_34(wires[202], wires[203], wires[176], wires[178], wires[114]);
full_adder fa_35(wires[204], wires[205], wires[175], wires[177], wires[179]);
full_adder fa_36(wires[206], wires[207], wires[180], wires[182], wires[184]);
full_adder fa_37(wires[208], wires[209], wires[181], wires[183], wires[185]);
full_adder fa_38(wires[210], wires[211], wires[186], wires[188], wires[160]);
full_adder fa_39(wires[212], wires[213], wires[187], wires[189], wires[190]);
full_adder fa_40(wires[214], wires[215], wires[191], wires[193], wires[194]);
full_adder fa_41(wires[216], wires[217], wires[197], wires[198], wires[136]);
full_adder fa_42(wires[218], wires[219], wires[199], wires[200], wires[202]);
full_adder fa_43(wires[220], wires[221], wires[201], wires[203], wires[204]);
full_adder fa_44(wires[222], wires[223], wires[205], wires[207], wires[208]);
full_adder fa_45(wires[224], wires[225], wires[209], wires[211], wires[212]);
half_adder ha_6(wires[226], wires[227], wires[213], wires[214]);
half_adder ha_7(wires[228], wires[229], wires[215], wires[195]);
half_adder ha_8(wires[230], wires[231], wires[217], wires[218]);
full_adder fa_46(wires[232], wires[233], wires[219], wires[220], wires[206]);
full_adder fa_47(wires[234], wires[235], wires[221], wires[222], wires[210]);
full_adder fa_48(wires[236], wires[237], wires[223], wires[224], wires[192]);
half_adder ha_9(wires[238], wires[239], wires[225], wires[226]);
half_adder ha_10(wires[240], wires[241], wires[227], wires[228]);
half_adder ha_11(wires[242], wires[243], wires[229], 1'b1);
half_adder ha_12(wires[244], wires[245], wires[231], wires[232]);
full_adder fa_49(wires[246], wires[247], wires[233], wires[234], wires[245]);
full_adder fa_50(wires[248], wires[249], wires[235], wires[236], wires[247]);
full_adder fa_51(wires[250], wires[251], wires[237], wires[238], wires[249]);
full_adder fa_52(wires[252], wires[253], wires[239], wires[240], wires[251]);
full_adder fa_53(wires[254], wires[255], wires[241], wires[242], wires[253]);
half_adder ha_13(wires[256], wires[257], wires[243], wires[255]);
endmodule