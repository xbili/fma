module pprt_16x16(out_0, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7);
input [15:0] in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7;
output [18:0] out_0;
wire [383:0] wires;
assign wires[0] = in_0[0];
assign wires[1] = in_0[1];
assign wires[2] = in_0[2];
assign wires[3] = in_0[3];
assign wires[4] = in_0[4];
assign wires[5] = in_0[5];
assign wires[6] = in_0[6];
assign wires[7] = in_0[7];
assign wires[8] = in_0[8];
assign wires[9] = in_0[9];
assign wires[10] = in_0[10];
assign wires[11] = in_0[11];
assign wires[12] = in_0[12];
assign wires[13] = in_0[13];
assign wires[14] = in_0[14];
assign wires[15] = in_0[15];
assign wires[16] = in_1[0];
assign wires[17] = in_1[1];
assign wires[18] = in_1[2];
assign wires[19] = in_1[3];
assign wires[20] = in_1[4];
assign wires[21] = in_1[5];
assign wires[22] = in_1[6];
assign wires[23] = in_1[7];
assign wires[24] = in_1[8];
assign wires[25] = in_1[9];
assign wires[26] = in_1[10];
assign wires[27] = in_1[11];
assign wires[28] = in_1[12];
assign wires[29] = in_1[13];
assign wires[30] = in_1[14];
assign wires[31] = in_1[15];
assign wires[32] = in_2[0];
assign wires[33] = in_2[1];
assign wires[34] = in_2[2];
assign wires[35] = in_2[3];
assign wires[36] = in_2[4];
assign wires[37] = in_2[5];
assign wires[38] = in_2[6];
assign wires[39] = in_2[7];
assign wires[40] = in_2[8];
assign wires[41] = in_2[9];
assign wires[42] = in_2[10];
assign wires[43] = in_2[11];
assign wires[44] = in_2[12];
assign wires[45] = in_2[13];
assign wires[46] = in_2[14];
assign wires[47] = in_2[15];
assign wires[48] = in_3[0];
assign wires[49] = in_3[1];
assign wires[50] = in_3[2];
assign wires[51] = in_3[3];
assign wires[52] = in_3[4];
assign wires[53] = in_3[5];
assign wires[54] = in_3[6];
assign wires[55] = in_3[7];
assign wires[56] = in_3[8];
assign wires[57] = in_3[9];
assign wires[58] = in_3[10];
assign wires[59] = in_3[11];
assign wires[60] = in_3[12];
assign wires[61] = in_3[13];
assign wires[62] = in_3[14];
assign wires[63] = in_3[15];
assign wires[64] = in_4[0];
assign wires[65] = in_4[1];
assign wires[66] = in_4[2];
assign wires[67] = in_4[3];
assign wires[68] = in_4[4];
assign wires[69] = in_4[5];
assign wires[70] = in_4[6];
assign wires[71] = in_4[7];
assign wires[72] = in_4[8];
assign wires[73] = in_4[9];
assign wires[74] = in_4[10];
assign wires[75] = in_4[11];
assign wires[76] = in_4[12];
assign wires[77] = in_4[13];
assign wires[78] = in_4[14];
assign wires[79] = in_4[15];
assign wires[80] = in_5[0];
assign wires[81] = in_5[1];
assign wires[82] = in_5[2];
assign wires[83] = in_5[3];
assign wires[84] = in_5[4];
assign wires[85] = in_5[5];
assign wires[86] = in_5[6];
assign wires[87] = in_5[7];
assign wires[88] = in_5[8];
assign wires[89] = in_5[9];
assign wires[90] = in_5[10];
assign wires[91] = in_5[11];
assign wires[92] = in_5[12];
assign wires[93] = in_5[13];
assign wires[94] = in_5[14];
assign wires[95] = in_5[15];
assign wires[96] = in_6[0];
assign wires[97] = in_6[1];
assign wires[98] = in_6[2];
assign wires[99] = in_6[3];
assign wires[100] = in_6[4];
assign wires[101] = in_6[5];
assign wires[102] = in_6[6];
assign wires[103] = in_6[7];
assign wires[104] = in_6[8];
assign wires[105] = in_6[9];
assign wires[106] = in_6[10];
assign wires[107] = in_6[11];
assign wires[108] = in_6[12];
assign wires[109] = in_6[13];
assign wires[110] = in_6[14];
assign wires[111] = in_6[15];
assign wires[112] = in_7[0];
assign wires[113] = in_7[1];
assign wires[114] = in_7[2];
assign wires[115] = in_7[3];
assign wires[116] = in_7[4];
assign wires[117] = in_7[5];
assign wires[118] = in_7[6];
assign wires[119] = in_7[7];
assign wires[120] = in_7[8];
assign wires[121] = in_7[9];
assign wires[122] = in_7[10];
assign wires[123] = in_7[11];
assign wires[124] = in_7[12];
assign wires[125] = in_7[13];
assign wires[126] = in_7[14];
assign wires[127] = in_7[15];
assign out_0[0] = wires[224];
assign out_0[1] = wires[288];
assign out_0[2] = wires[320];
assign out_0[3] = wires[352];
assign out_0[4] = wires[354];
assign out_0[5] = wires[356];
assign out_0[6] = wires[358];
assign out_0[7] = wires[360];
assign out_0[8] = wires[362];
assign out_0[9] = wires[364];
assign out_0[10] = wires[366];
assign out_0[11] = wires[368];
assign out_0[12] = wires[370];
assign out_0[13] = wires[372];
assign out_0[14] = wires[374];
assign out_0[15] = wires[376];
assign out_0[16] = wires[378];
assign out_0[17] = wires[380];
assign out_0[18] = wires[382];
full_adder fa_0(wires[128], wires[129], wires[0], wires[16], wires[32]);
full_adder fa_1(wires[130], wires[131], wires[48], wires[64], wires[80]);
half_adder ha_0(wires[132], wires[133], wires[96], wires[112]);
full_adder fa_2(wires[134], wires[135], wires[1], wires[17], wires[33]);
full_adder fa_3(wires[136], wires[137], wires[49], wires[65], wires[81]);
half_adder ha_1(wires[138], wires[139], wires[97], wires[113]);
full_adder fa_4(wires[140], wires[141], wires[2], wires[18], wires[34]);
full_adder fa_5(wires[142], wires[143], wires[50], wires[66], wires[82]);
half_adder ha_2(wires[144], wires[145], wires[98], wires[114]);
full_adder fa_6(wires[146], wires[147], wires[3], wires[19], wires[35]);
full_adder fa_7(wires[148], wires[149], wires[51], wires[67], wires[83]);
half_adder ha_3(wires[150], wires[151], wires[99], wires[115]);
full_adder fa_8(wires[152], wires[153], wires[4], wires[20], wires[36]);
full_adder fa_9(wires[154], wires[155], wires[52], wires[68], wires[84]);
half_adder ha_4(wires[156], wires[157], wires[100], wires[116]);
full_adder fa_10(wires[158], wires[159], wires[5], wires[21], wires[37]);
full_adder fa_11(wires[160], wires[161], wires[53], wires[69], wires[85]);
half_adder ha_5(wires[162], wires[163], wires[101], wires[117]);
full_adder fa_12(wires[164], wires[165], wires[6], wires[22], wires[38]);
full_adder fa_13(wires[166], wires[167], wires[54], wires[70], wires[86]);
half_adder ha_6(wires[168], wires[169], wires[102], wires[118]);
full_adder fa_14(wires[170], wires[171], wires[7], wires[23], wires[39]);
full_adder fa_15(wires[172], wires[173], wires[55], wires[71], wires[87]);
half_adder ha_7(wires[174], wires[175], wires[103], wires[119]);
full_adder fa_16(wires[176], wires[177], wires[8], wires[24], wires[40]);
full_adder fa_17(wires[178], wires[179], wires[56], wires[72], wires[88]);
half_adder ha_8(wires[180], wires[181], wires[104], wires[120]);
full_adder fa_18(wires[182], wires[183], wires[9], wires[25], wires[41]);
full_adder fa_19(wires[184], wires[185], wires[57], wires[73], wires[89]);
half_adder ha_9(wires[186], wires[187], wires[105], wires[121]);
full_adder fa_20(wires[188], wires[189], wires[10], wires[26], wires[42]);
full_adder fa_21(wires[190], wires[191], wires[58], wires[74], wires[90]);
half_adder ha_10(wires[192], wires[193], wires[106], wires[122]);
full_adder fa_22(wires[194], wires[195], wires[11], wires[27], wires[43]);
full_adder fa_23(wires[196], wires[197], wires[59], wires[75], wires[91]);
half_adder ha_11(wires[198], wires[199], wires[107], wires[123]);
full_adder fa_24(wires[200], wires[201], wires[12], wires[28], wires[44]);
full_adder fa_25(wires[202], wires[203], wires[60], wires[76], wires[92]);
half_adder ha_12(wires[204], wires[205], wires[108], wires[124]);
full_adder fa_26(wires[206], wires[207], wires[13], wires[29], wires[45]);
full_adder fa_27(wires[208], wires[209], wires[61], wires[77], wires[93]);
half_adder ha_13(wires[210], wires[211], wires[109], wires[125]);
full_adder fa_28(wires[212], wires[213], wires[14], wires[30], wires[46]);
full_adder fa_29(wires[214], wires[215], wires[62], wires[78], wires[94]);
half_adder ha_14(wires[216], wires[217], wires[110], wires[126]);
full_adder fa_30(wires[218], wires[219], wires[15], wires[31], wires[47]);
full_adder fa_31(wires[220], wires[221], wires[63], wires[79], wires[95]);
half_adder ha_15(wires[222], wires[223], wires[111], wires[127]);
full_adder fa_32(wires[224], wires[225], wires[128], wires[130], wires[132]);
full_adder fa_33(wires[226], wires[227], wires[129], wires[131], wires[133]);
full_adder fa_34(wires[228], wires[229], wires[134], wires[136], wires[138]);
full_adder fa_35(wires[230], wires[231], wires[135], wires[137], wires[139]);
full_adder fa_36(wires[232], wires[233], wires[140], wires[142], wires[144]);
full_adder fa_37(wires[234], wires[235], wires[141], wires[143], wires[145]);
full_adder fa_38(wires[236], wires[237], wires[146], wires[148], wires[150]);
full_adder fa_39(wires[238], wires[239], wires[147], wires[149], wires[151]);
full_adder fa_40(wires[240], wires[241], wires[152], wires[154], wires[156]);
full_adder fa_41(wires[242], wires[243], wires[153], wires[155], wires[157]);
full_adder fa_42(wires[244], wires[245], wires[158], wires[160], wires[162]);
full_adder fa_43(wires[246], wires[247], wires[159], wires[161], wires[163]);
full_adder fa_44(wires[248], wires[249], wires[164], wires[166], wires[168]);
full_adder fa_45(wires[250], wires[251], wires[165], wires[167], wires[169]);
full_adder fa_46(wires[252], wires[253], wires[170], wires[172], wires[174]);
full_adder fa_47(wires[254], wires[255], wires[171], wires[173], wires[175]);
full_adder fa_48(wires[256], wires[257], wires[176], wires[178], wires[180]);
full_adder fa_49(wires[258], wires[259], wires[177], wires[179], wires[181]);
full_adder fa_50(wires[260], wires[261], wires[182], wires[184], wires[186]);
full_adder fa_51(wires[262], wires[263], wires[183], wires[185], wires[187]);
full_adder fa_52(wires[264], wires[265], wires[188], wires[190], wires[192]);
full_adder fa_53(wires[266], wires[267], wires[189], wires[191], wires[193]);
full_adder fa_54(wires[268], wires[269], wires[194], wires[196], wires[198]);
full_adder fa_55(wires[270], wires[271], wires[195], wires[197], wires[199]);
full_adder fa_56(wires[272], wires[273], wires[200], wires[202], wires[204]);
full_adder fa_57(wires[274], wires[275], wires[201], wires[203], wires[205]);
full_adder fa_58(wires[276], wires[277], wires[206], wires[208], wires[210]);
full_adder fa_59(wires[278], wires[279], wires[207], wires[209], wires[211]);
full_adder fa_60(wires[280], wires[281], wires[212], wires[214], wires[216]);
full_adder fa_61(wires[282], wires[283], wires[213], wires[215], wires[217]);
full_adder fa_62(wires[284], wires[285], wires[218], wires[220], wires[222]);
full_adder fa_63(wires[286], wires[287], wires[219], wires[221], wires[223]);
full_adder fa_64(wires[288], wires[289], wires[225], wires[226], wires[228]);
full_adder fa_65(wires[290], wires[291], wires[227], wires[229], wires[230]);
full_adder fa_66(wires[292], wires[293], wires[231], wires[233], wires[234]);
full_adder fa_67(wires[294], wires[295], wires[235], wires[237], wires[238]);
full_adder fa_68(wires[296], wires[297], wires[239], wires[241], wires[242]);
full_adder fa_69(wires[298], wires[299], wires[243], wires[245], wires[246]);
full_adder fa_70(wires[300], wires[301], wires[247], wires[249], wires[250]);
full_adder fa_71(wires[302], wires[303], wires[251], wires[253], wires[254]);
full_adder fa_72(wires[304], wires[305], wires[255], wires[257], wires[258]);
full_adder fa_73(wires[306], wires[307], wires[259], wires[261], wires[262]);
full_adder fa_74(wires[308], wires[309], wires[263], wires[265], wires[266]);
full_adder fa_75(wires[310], wires[311], wires[267], wires[269], wires[270]);
full_adder fa_76(wires[312], wires[313], wires[271], wires[273], wires[274]);
full_adder fa_77(wires[314], wires[315], wires[275], wires[277], wires[278]);
full_adder fa_78(wires[316], wires[317], wires[279], wires[281], wires[282]);
full_adder fa_79(wires[318], wires[319], wires[283], wires[285], wires[286]);
full_adder fa_80(wires[320], wires[321], wires[289], wires[290], wires[232]);
full_adder fa_81(wires[322], wires[323], wires[291], wires[292], wires[236]);
full_adder fa_82(wires[324], wires[325], wires[293], wires[294], wires[240]);
full_adder fa_83(wires[326], wires[327], wires[295], wires[296], wires[244]);
full_adder fa_84(wires[328], wires[329], wires[297], wires[298], wires[248]);
full_adder fa_85(wires[330], wires[331], wires[299], wires[300], wires[252]);
full_adder fa_86(wires[332], wires[333], wires[301], wires[302], wires[256]);
full_adder fa_87(wires[334], wires[335], wires[303], wires[304], wires[260]);
full_adder fa_88(wires[336], wires[337], wires[305], wires[306], wires[264]);
full_adder fa_89(wires[338], wires[339], wires[307], wires[308], wires[268]);
full_adder fa_90(wires[340], wires[341], wires[309], wires[310], wires[272]);
full_adder fa_91(wires[342], wires[343], wires[311], wires[312], wires[276]);
full_adder fa_92(wires[344], wires[345], wires[313], wires[314], wires[280]);
full_adder fa_93(wires[346], wires[347], wires[315], wires[316], wires[284]);
half_adder ha_16(wires[348], wires[349], wires[317], wires[318]);
half_adder ha_17(wires[350], wires[351], wires[319], wires[287]);
half_adder ha_18(wires[352], wires[353], wires[321], wires[322]);
full_adder fa_94(wires[354], wires[355], wires[323], wires[324], wires[353]);
full_adder fa_95(wires[356], wires[357], wires[325], wires[326], wires[355]);
full_adder fa_96(wires[358], wires[359], wires[327], wires[328], wires[357]);
full_adder fa_97(wires[360], wires[361], wires[329], wires[330], wires[359]);
full_adder fa_98(wires[362], wires[363], wires[331], wires[332], wires[361]);
full_adder fa_99(wires[364], wires[365], wires[333], wires[334], wires[363]);
full_adder fa_100(wires[366], wires[367], wires[335], wires[336], wires[365]);
full_adder fa_101(wires[368], wires[369], wires[337], wires[338], wires[367]);
full_adder fa_102(wires[370], wires[371], wires[339], wires[340], wires[369]);
full_adder fa_103(wires[372], wires[373], wires[341], wires[342], wires[371]);
full_adder fa_104(wires[374], wires[375], wires[343], wires[344], wires[373]);
full_adder fa_105(wires[376], wires[377], wires[345], wires[346], wires[375]);
full_adder fa_106(wires[378], wires[379], wires[347], wires[348], wires[377]);
full_adder fa_107(wires[380], wires[381], wires[349], wires[350], wires[379]);
half_adder ha_19(wires[382], wires[383], wires[351], wires[381]);
endmodule